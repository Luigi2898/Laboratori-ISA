library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;
    use work.array_std.all;


entity DADDA is
  generic(N : integer := 32; N_PP : integer := 17);
  port (
    PP1      : in  std_logic_vector (N downto 0);
    PP2      : in  std_logic_vector (N downto 0);
    PP3      : in  std_logic_vector (N downto 0);
    PP4      : in  std_logic_vector (N downto 0);
    PP5      : in  std_logic_vector (N downto 0);
    PP6      : in  std_logic_vector (N downto 0);
    PP7      : in  std_logic_vector (N downto 0);
    PP8      : in  std_logic_vector (N downto 0);
    PP9      : in  std_logic_vector (N downto 0);
    PP10     : in  std_logic_vector (N downto 0);
    PP11     : in  std_logic_vector (N downto 0);
    PP12     : in  std_logic_vector (N downto 0);
    PP13     : in  std_logic_vector (N downto 0);
    PP14     : in  std_logic_vector (N downto 0);
    PP15     : in  std_logic_vector (N downto 0);
    PP16     : in  std_logic_vector (N downto 0);
    PP17     : in  std_logic_vector (N downto 0);
    PP_sign : in  std_logic_vector (N / 2 downto 0);
    SUM     : out std_logic_vector (2 * N - 1 downto 0)
  ) ;
end DADDA;

architecture structural of DADDA is
  
  component FA IS
    port(
		A, B, Cin : IN STD_LOGIC;
		S, Co : OUT STD_LOGIC
	);	
  end component FA;

  component HA is
    port(
		    A, B  : in  std_logic;
		    S, Co : out std_logic
    );
  end component HA;
signal internal_0_0 : std_logic_vector(64 downto 0);
signal internal_0_1 : std_logic_vector(64 downto 0);
signal internal_0_2 : std_logic_vector(64 downto 0);
signal internal_0_3 : std_logic_vector(64 downto 0);
signal internal_0_4 : std_logic_vector(64 downto 0);
signal internal_0_5 : std_logic_vector(64 downto 0);
signal internal_0_6 : std_logic_vector(64 downto 0);
signal internal_0_7 : std_logic_vector(64 downto 0);
signal internal_0_8 : std_logic_vector(64 downto 0);
signal internal_0_9 : std_logic_vector(64 downto 0);
signal internal_0_10 : std_logic_vector(64 downto 0);
signal internal_0_11 : std_logic_vector(64 downto 0);
signal internal_0_12 : std_logic_vector(64 downto 0);
signal internal_0_13 : std_logic_vector(64 downto 0);
signal internal_0_14 : std_logic_vector(64 downto 0);
signal internal_0_15 : std_logic_vector(64 downto 0);
signal internal_0_16 : std_logic_vector(64 downto 0);
signal internal_1_0 : std_logic_vector(64 downto 0);
signal internal_1_1 : std_logic_vector(64 downto 0);
signal internal_1_2 : std_logic_vector(64 downto 0);
signal internal_1_3 : std_logic_vector(64 downto 0);
signal internal_1_4 : std_logic_vector(64 downto 0);
signal internal_1_5 : std_logic_vector(64 downto 0);
signal internal_1_6 : std_logic_vector(64 downto 0);
signal internal_1_7 : std_logic_vector(64 downto 0);
signal internal_1_8 : std_logic_vector(64 downto 0);
signal internal_1_9 : std_logic_vector(64 downto 0);
signal internal_1_10 : std_logic_vector(64 downto 0);
signal internal_1_11 : std_logic_vector(64 downto 0);
signal internal_1_12 : std_logic_vector(64 downto 0);
signal internal_2_0 : std_logic_vector(64 downto 0);
signal internal_2_1 : std_logic_vector(64 downto 0);
signal internal_2_2 : std_logic_vector(64 downto 0);
signal internal_2_3 : std_logic_vector(64 downto 0);
signal internal_2_4 : std_logic_vector(64 downto 0);
signal internal_2_5 : std_logic_vector(64 downto 0);
signal internal_2_6 : std_logic_vector(64 downto 0);
signal internal_2_7 : std_logic_vector(64 downto 0);
signal internal_2_8 : std_logic_vector(64 downto 0);
signal internal_3_0 : std_logic_vector(64 downto 0);
signal internal_3_1 : std_logic_vector(64 downto 0);
signal internal_3_2 : std_logic_vector(64 downto 0);
signal internal_3_3 : std_logic_vector(64 downto 0);
signal internal_3_4 : std_logic_vector(64 downto 0);
signal internal_3_5 : std_logic_vector(64 downto 0);
signal internal_4_0 : std_logic_vector(64 downto 0);
signal internal_4_1 : std_logic_vector(64 downto 0);
signal internal_4_2 : std_logic_vector(64 downto 0);
signal internal_4_3 : std_logic_vector(64 downto 0);
signal internal_5_0 : std_logic_vector(64 downto 0);
signal internal_5_1 : std_logic_vector(64 downto 0);
signal internal_5_2 : std_logic_vector(64 downto 0);
signal internal_6_0 : std_logic_vector(64 downto 0);
signal internal_6_1 : std_logic_vector(64 downto 0);




begin

internal_0_0 <= '0' & not(PP_sign(15)) & '1' & not(PP_sign(14)) & '1' & not(PP_sign(13)) & '1' & not(PP_sign(12)) & '1' & not(PP_sign(11)) & '1' & not(PP_sign(10)) & '1' & not(PP_sign(9)) & '1' & not(PP_sign(8)) & '1' & not(PP_sign(7)) & '1' & not(PP_sign(6)) & '1' & not(PP_sign(5)) & '1' & not(PP_sign(4)) & '1' & not(PP_sign(3)) & '1' & not(PP_sign(2)) & '1' & not(PP_sign(0)) & PP_sign(0) & PP_sign(0) & PP1(32) & PP1(31) & PP1(30) & PP1(29) & PP1(28) & PP1(27) & PP1(26) & PP1(25) & PP1(24) & PP1(23) & PP1(22) & PP1(21) & PP1(20) & PP1(19) & PP1(18) & PP1(17) & PP1(16) & PP1(15) & PP1(14) & PP1(13) & PP1(12) & PP1(11) & PP1(10) & PP1(9) & PP1(8) & PP1(7) & PP1(6) & PP1(5) & PP1(4) & PP1(3) & PP1(2) & PP1(1) & PP1(0) ;
internal_0_1 <= '0' & PP17(31) & PP16(32) & PP16(31) & PP15(32) & PP15(31) & PP14(32) & PP14(31) & PP13(32) & PP13(31) & PP12(32) & PP12(31) & PP11(32) & PP11(31) & PP10(32) & PP10(31) & PP9(32) & PP9(31) & PP8(32) & PP8(31) & PP7(32) & PP7(31) & PP6(32) & PP6(31) & PP5(32) & PP5(31) & PP4(32) & PP4(31) & PP3(32) & not(PP_sign(1)) & PP2(32) & PP2(31) & PP2(30) & PP2(29) & PP2(28) & PP2(27) & PP2(26) & PP2(25) & PP2(24) & PP2(23) & PP2(22) & PP2(21) & PP2(20) & PP2(19) & PP2(18) & PP2(17) & PP2(16) & PP2(15) & PP2(14) & PP2(13) & PP2(12) & PP2(11) & PP2(10) & PP2(9) & PP2(8) & PP2(7) & PP2(6) & PP2(5) & PP2(4) & PP2(3) & PP2(2) & PP2(1) & PP2(0) & '0' & PP_sign(0) ;
internal_0_2 <= '0' & '0' & PP17(30) & PP17(29) & PP16(30) & PP16(29) & PP15(30) & PP15(29) & PP14(30) & PP14(29) & PP13(30) & PP13(29) & PP12(30) & PP12(29) & PP11(30) & PP11(29) & PP10(30) & PP10(29) & PP9(30) & PP9(29) & PP8(30) & PP8(29) & PP7(30) & PP7(29) & PP6(30) & PP6(29) & PP5(30) & PP5(29) & PP4(30) & PP3(31) & PP3(30) & PP3(29) & PP3(28) & PP3(27) & PP3(26) & PP3(25) & PP3(24) & PP3(23) & PP3(22) & PP3(21) & PP3(20) & PP3(19) & PP3(18) & PP3(17) & PP3(16) & PP3(15) & PP3(14) & PP3(13) & PP3(12) & PP3(11) & PP3(10) & PP3(9) & PP3(8) & PP3(7) & PP3(6) & PP3(5) & PP3(4) & PP3(3) & PP3(2) & PP3(1) & PP3(0) & '0' & PP_sign(1) & '0' & '0' ;
internal_0_3 <= '0' & '0' & '0' & '0' & PP17(28) & PP17(27) & PP16(28) & PP16(27) & PP15(28) & PP15(27) & PP14(28) & PP14(27) & PP13(28) & PP13(27) & PP12(28) & PP12(27) & PP11(28) & PP11(27) & PP10(28) & PP10(27) & PP9(28) & PP9(27) & PP8(28) & PP8(27) & PP7(28) & PP7(27) & PP6(28) & PP6(27) & PP5(28) & PP4(29) & PP4(28) & PP4(27) & PP4(26) & PP4(25) & PP4(24) & PP4(23) & PP4(22) & PP4(21) & PP4(20) & PP4(19) & PP4(18) & PP4(17) & PP4(16) & PP4(15) & PP4(14) & PP4(13) & PP4(12) & PP4(11) & PP4(10) & PP4(9) & PP4(8) & PP4(7) & PP4(6) & PP4(5) & PP4(4) & PP4(3) & PP4(2) & PP4(1) & PP4(0) & '0' & PP_sign(2) & '0' & '0' & '0' & '0' ;
internal_0_4 <= '0' & '0' & '0' & '0' & '0' & '0' & PP17(26) & PP17(25) & PP16(26) & PP16(25) & PP15(26) & PP15(25) & PP14(26) & PP14(25) & PP13(26) & PP13(25) & PP12(26) & PP12(25) & PP11(26) & PP11(25) & PP10(26) & PP10(25) & PP9(26) & PP9(25) & PP8(26) & PP8(25) & PP7(26) & PP7(25) & PP6(26) & PP5(27) & PP5(26) & PP5(25) & PP5(24) & PP5(23) & PP5(22) & PP5(21) & PP5(20) & PP5(19) & PP5(18) & PP5(17) & PP5(16) & PP5(15) & PP5(14) & PP5(13) & PP5(12) & PP5(11) & PP5(10) & PP5(9) & PP5(8) & PP5(7) & PP5(6) & PP5(5) & PP5(4) & PP5(3) & PP5(2) & PP5(1) & PP5(0) & '0' & PP_sign(3) & '0' & '0' & '0' & '0' & '0' & '0' ;
internal_0_5 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & PP17(24) & PP17(23) & PP16(24) & PP16(23) & PP15(24) & PP15(23) & PP14(24) & PP14(23) & PP13(24) & PP13(23) & PP12(24) & PP12(23) & PP11(24) & PP11(23) & PP10(24) & PP10(23) & PP9(24) & PP9(23) & PP8(24) & PP8(23) & PP7(24) & PP6(25) & PP6(24) & PP6(23) & PP6(22) & PP6(21) & PP6(20) & PP6(19) & PP6(18) & PP6(17) & PP6(16) & PP6(15) & PP6(14) & PP6(13) & PP6(12) & PP6(11) & PP6(10) & PP6(9) & PP6(8) & PP6(7) & PP6(6) & PP6(5) & PP6(4) & PP6(3) & PP6(2) & PP6(1) & PP6(0) & '0' & PP_sign(4) & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' ;
internal_0_6 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & PP17(22) & PP17(21) & PP16(22) & PP16(21) & PP15(22) & PP15(21) & PP14(22) & PP14(21) & PP13(22) & PP13(21) & PP12(22) & PP12(21) & PP11(22) & PP11(21) & PP10(22) & PP10(21) & PP9(22) & PP9(21) & PP8(22) & PP7(23) & PP7(22) & PP7(21) & PP7(20) & PP7(19) & PP7(18) & PP7(17) & PP7(16) & PP7(15) & PP7(14) & PP7(13) & PP7(12) & PP7(11) & PP7(10) & PP7(9) & PP7(8) & PP7(7) & PP7(6) & PP7(5) & PP7(4) & PP7(3) & PP7(2) & PP7(1) & PP7(0) & '0' & PP_sign(5) & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' ;
internal_0_7 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & PP17(20) & PP17(19) & PP16(20) & PP16(19) & PP15(20) & PP15(19) & PP14(20) & PP14(19) & PP13(20) & PP13(19) & PP12(20) & PP12(19) & PP11(20) & PP11(19) & PP10(20) & PP10(19) & PP9(20) & PP8(21) & PP8(20) & PP8(19) & PP8(18) & PP8(17) & PP8(16) & PP8(15) & PP8(14) & PP8(13) & PP8(12) & PP8(11) & PP8(10) & PP8(9) & PP8(8) & PP8(7) & PP8(6) & PP8(5) & PP8(4) & PP8(3) & PP8(2) & PP8(1) & PP8(0) & '0' & PP_sign(6) & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' ;
internal_0_8 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & PP17(18) & PP17(17) & PP16(18) & PP16(17) & PP15(18) & PP15(17) & PP14(18) & PP14(17) & PP13(18) & PP13(17) & PP12(18) & PP12(17) & PP11(18) & PP11(17) & PP10(18) & PP9(19) & PP9(18) & PP9(17) & PP9(16) & PP9(15) & PP9(14) & PP9(13) & PP9(12) & PP9(11) & PP9(10) & PP9(9) & PP9(8) & PP9(7) & PP9(6) & PP9(5) & PP9(4) & PP9(3) & PP9(2) & PP9(1) & PP9(0) & '0' & PP_sign(7) & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' ;
internal_0_9 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & PP17(16) & PP17(15) & PP16(16) & PP16(15) & PP15(16) & PP15(15) & PP14(16) & PP14(15) & PP13(16) & PP13(15) & PP12(16) & PP12(15) & PP11(16) & PP10(17) & PP10(16) & PP10(15) & PP10(14) & PP10(13) & PP10(12) & PP10(11) & PP10(10) & PP10(9) & PP10(8) & PP10(7) & PP10(6) & PP10(5) & PP10(4) & PP10(3) & PP10(2) & PP10(1) & PP10(0) & '0' & PP_sign(8) & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' ;
internal_0_10 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & PP17(14) & PP17(13) & PP16(14) & PP16(13) & PP15(14) & PP15(13) & PP14(14) & PP14(13) & PP13(14) & PP13(13) & PP12(14) & PP11(15) & PP11(14) & PP11(13) & PP11(12) & PP11(11) & PP11(10) & PP11(9) & PP11(8) & PP11(7) & PP11(6) & PP11(5) & PP11(4) & PP11(3) & PP11(2) & PP11(1) & PP11(0) & '0' & PP_sign(9) & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' ;
internal_0_11 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & PP17(12) & PP17(11) & PP16(12) & PP16(11) & PP15(12) & PP15(11) & PP14(12) & PP14(11) & PP13(12) & PP12(13) & PP12(12) & PP12(11) & PP12(10) & PP12(9) & PP12(8) & PP12(7) & PP12(6) & PP12(5) & PP12(4) & PP12(3) & PP12(2) & PP12(1) & PP12(0) & '0' & PP_sign(10) & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' ;
internal_0_12 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & PP17(10) & PP17(9) & PP16(10) & PP16(9) & PP15(10) & PP15(9) & PP14(10) & PP13(11) & PP13(10) & PP13(9) & PP13(8) & PP13(7) & PP13(6) & PP13(5) & PP13(4) & PP13(3) & PP13(2) & PP13(1) & PP13(0) & '0' & PP_sign(11) & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' ;
internal_0_13 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & PP17(8) & PP17(7) & PP16(8) & PP16(7) & PP15(8) & PP14(9) & PP14(8) & PP14(7) & PP14(6) & PP14(5) & PP14(4) & PP14(3) & PP14(2) & PP14(1) & PP14(0) & '0' & PP_sign(12) & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' ;
internal_0_14 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & PP17(6) & PP17(5) & PP16(6) & PP15(7) & PP15(6) & PP15(5) & PP15(4) & PP15(3) & PP15(2) & PP15(1) & PP15(0) & '0' & PP_sign(13) & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' ;
internal_0_15 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & PP17(4) & PP16(5) & PP16(4) & PP16(3) & PP16(2) & PP16(1) & PP16(0) & '0' & PP_sign(14) & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' ;
internal_0_16 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & PP17(3) & PP17(2) & PP17(1) & PP17(0) & '0' & PP_sign(15) & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' ;


HA_0 : HA port map(internal_0_0( 24 ), internal_0_1( 24 ), internal_1_0( 24 ), internal_1_1( 25 ));
HA_1 : HA port map(internal_0_0( 25 ), internal_0_1( 25 ), internal_1_0( 25 ), internal_1_1( 26 ));
FA_0 : FA port map(internal_0_0( 26 ), internal_0_1( 26 ), internal_0_2( 26 ), internal_1_0( 26 ), internal_1_1( 27 ));
HA_2 : HA port map(internal_0_3( 26 ), internal_0_4( 26 ), internal_1_1( 26 ), internal_1_2( 27 ));
FA_1 : FA port map(internal_0_0( 27 ), internal_0_1( 27 ), internal_0_2( 27 ), internal_1_0( 27 ), internal_1_1( 28 ));
HA_3 : HA port map(internal_0_3( 27 ), internal_0_4( 27 ), internal_1_1( 27 ), internal_1_2( 28 ));
FA_2 : FA port map(internal_0_0( 28 ), internal_0_1( 28 ), internal_0_2( 28 ), internal_1_0( 28 ), internal_1_1( 29 ));
FA_3 : FA port map(internal_0_3( 28 ), internal_0_4( 28 ), internal_0_5( 28 ), internal_1_0( 28 ), internal_1_1( 29 ));
HA_4 : HA port map(internal_0_6( 28 ), internal_0_7( 28 ), internal_1_2( 28 ), internal_1_3( 29 ));
FA_4 : FA port map(internal_0_0( 29 ), internal_0_1( 29 ), internal_0_2( 29 ), internal_1_0( 29 ), internal_1_1( 30 ));
FA_5 : FA port map(internal_0_3( 29 ), internal_0_4( 29 ), internal_0_5( 29 ), internal_1_0( 29 ), internal_1_1( 30 ));
HA_5 : HA port map(internal_0_6( 29 ), internal_0_7( 29 ), internal_1_2( 29 ), internal_1_3( 30 ));
FA_6 : FA port map(internal_0_0( 30 ), internal_0_1( 30 ), internal_0_2( 30 ), internal_1_0( 30 ), internal_1_1( 31 ));
FA_7 : FA port map(internal_0_3( 30 ), internal_0_4( 30 ), internal_0_5( 30 ), internal_1_0( 30 ), internal_1_1( 31 ));
FA_8 : FA port map(internal_0_6( 30 ), internal_0_7( 30 ), internal_0_8( 30 ), internal_1_0( 30 ), internal_1_1( 31 ));
HA_6 : HA port map(internal_0_9( 30 ), internal_0_10( 30 ), internal_1_3( 30 ), internal_1_4( 31 ));
FA_9 : FA port map(internal_0_0( 31 ), internal_0_1( 31 ), internal_0_2( 31 ), internal_1_0( 31 ), internal_1_1( 32 ));
FA_10 : FA port map(internal_0_3( 31 ), internal_0_4( 31 ), internal_0_5( 31 ), internal_1_0( 31 ), internal_1_1( 32 ));
FA_11 : FA port map(internal_0_6( 31 ), internal_0_7( 31 ), internal_0_8( 31 ), internal_1_0( 31 ), internal_1_1( 32 ));
HA_7 : HA port map(internal_0_9( 31 ), internal_0_10( 31 ), internal_1_3( 31 ), internal_1_4( 32 ));
FA_12 : FA port map(internal_0_0( 32 ), internal_0_1( 32 ), internal_0_2( 32 ), internal_1_0( 32 ), internal_1_1( 33 ));
FA_13 : FA port map(internal_0_3( 32 ), internal_0_4( 32 ), internal_0_5( 32 ), internal_1_0( 32 ), internal_1_1( 33 ));
FA_14 : FA port map(internal_0_6( 32 ), internal_0_7( 32 ), internal_0_8( 32 ), internal_1_0( 32 ), internal_1_1( 33 ));
FA_15 : FA port map(internal_0_9( 32 ), internal_0_10( 32 ), internal_0_11( 32 ), internal_1_1( 32 ), internal_1_2( 33 ));
FA_16 : FA port map(internal_0_0( 33 ), internal_0_1( 33 ), internal_0_2( 33 ), internal_1_0( 33 ), internal_1_1( 34 ));
FA_17 : FA port map(internal_0_3( 33 ), internal_0_4( 33 ), internal_0_5( 33 ), internal_1_0( 33 ), internal_1_1( 34 ));
FA_18 : FA port map(internal_0_6( 33 ), internal_0_7( 33 ), internal_0_8( 33 ), internal_1_0( 33 ), internal_1_1( 34 ));
FA_19 : FA port map(internal_0_9( 33 ), internal_0_10( 33 ), internal_0_11( 33 ), internal_1_1( 33 ), internal_1_2( 34 ));
FA_20 : FA port map(internal_0_0( 34 ), internal_0_1( 34 ), internal_0_2( 34 ), internal_1_0( 34 ), internal_1_1( 35 ));
FA_21 : FA port map(internal_0_3( 34 ), internal_0_4( 34 ), internal_0_5( 34 ), internal_1_0( 34 ), internal_1_1( 35 ));
FA_22 : FA port map(internal_0_6( 34 ), internal_0_7( 34 ), internal_0_8( 34 ), internal_1_0( 34 ), internal_1_1( 35 ));
FA_23 : FA port map(internal_0_9( 34 ), internal_0_10( 34 ), internal_0_11( 34 ), internal_1_1( 34 ), internal_1_2( 35 ));
FA_24 : FA port map(internal_0_0( 35 ), internal_0_1( 35 ), internal_0_2( 35 ), internal_1_0( 35 ), internal_1_1( 36 ));
FA_25 : FA port map(internal_0_3( 35 ), internal_0_4( 35 ), internal_0_5( 35 ), internal_1_0( 35 ), internal_1_1( 36 ));
FA_26 : FA port map(internal_0_6( 35 ), internal_0_7( 35 ), internal_0_8( 35 ), internal_1_0( 35 ), internal_1_1( 36 ));
FA_27 : FA port map(internal_0_9( 35 ), internal_0_10( 35 ), internal_0_11( 35 ), internal_1_1( 35 ), internal_1_2( 36 ));
FA_28 : FA port map(internal_0_0( 36 ), internal_0_1( 36 ), internal_0_2( 36 ), internal_1_0( 36 ), internal_1_1( 37 ));
FA_29 : FA port map(internal_0_3( 36 ), internal_0_4( 36 ), internal_0_5( 36 ), internal_1_0( 36 ), internal_1_1( 37 ));
FA_30 : FA port map(internal_0_6( 36 ), internal_0_7( 36 ), internal_0_8( 36 ), internal_1_0( 36 ), internal_1_1( 37 ));
HA_8 : HA port map(internal_0_9( 36 ), internal_0_10( 36 ), internal_1_3( 36 ), internal_1_4( 37 ));
FA_31 : FA port map(internal_0_0( 37 ), internal_0_1( 37 ), internal_0_2( 37 ), internal_1_0( 37 ), internal_1_1( 38 ));
FA_32 : FA port map(internal_0_3( 37 ), internal_0_4( 37 ), internal_0_5( 37 ), internal_1_0( 37 ), internal_1_1( 38 ));
FA_33 : FA port map(internal_0_6( 37 ), internal_0_7( 37 ), internal_0_8( 37 ), internal_1_0( 37 ), internal_1_1( 38 ));
FA_34 : FA port map(internal_0_0( 38 ), internal_0_1( 38 ), internal_0_2( 38 ), internal_1_0( 38 ), internal_1_1( 39 ));
FA_35 : FA port map(internal_0_3( 38 ), internal_0_4( 38 ), internal_0_5( 38 ), internal_1_0( 38 ), internal_1_1( 39 ));
HA_9 : HA port map(internal_0_6( 38 ), internal_0_7( 38 ), internal_1_2( 38 ), internal_1_3( 39 ));
FA_36 : FA port map(internal_0_0( 39 ), internal_0_1( 39 ), internal_0_2( 39 ), internal_1_0( 39 ), internal_1_1( 40 ));
FA_37 : FA port map(internal_0_3( 39 ), internal_0_4( 39 ), internal_0_5( 39 ), internal_1_0( 39 ), internal_1_1( 40 ));
FA_38 : FA port map(internal_0_0( 40 ), internal_0_1( 40 ), internal_0_2( 40 ), internal_1_0( 40 ), internal_1_1( 41 ));
HA_10 : HA port map(internal_0_3( 40 ), internal_0_4( 40 ), internal_1_1( 40 ), internal_1_2( 41 ));
FA_39 : FA port map(internal_0_0( 41 ), internal_0_1( 41 ), internal_0_2( 41 ), internal_1_0( 41 ), internal_1_1( 42 ));
HA_11 : HA port map(internal_0_0( 42 ), internal_0_1( 42 ), internal_1_0( 42 ), internal_1_1( 43 ));
HA_12 : HA port map(internal_1_0( 16 ), internal_1_1( 16 ), internal_2_0( 16 ), internal_2_1( 17 ));
HA_13 : HA port map(internal_1_0( 17 ), internal_1_1( 17 ), internal_2_0( 17 ), internal_2_1( 18 ));
FA_40 : FA port map(internal_1_0( 18 ), internal_1_1( 18 ), internal_1_2( 18 ), internal_2_0( 18 ), internal_2_1( 19 ));
HA_14 : HA port map(internal_1_3( 18 ), internal_1_4( 18 ), internal_2_1( 18 ), internal_2_2( 19 ));
FA_41 : FA port map(internal_1_0( 19 ), internal_1_1( 19 ), internal_1_2( 19 ), internal_2_0( 19 ), internal_2_1( 20 ));
HA_15 : HA port map(internal_1_3( 19 ), internal_1_4( 19 ), internal_2_1( 19 ), internal_2_2( 20 ));
FA_42 : FA port map(internal_1_0( 20 ), internal_1_1( 20 ), internal_1_2( 20 ), internal_2_0( 20 ), internal_2_1( 21 ));
FA_43 : FA port map(internal_1_3( 20 ), internal_1_4( 20 ), internal_1_5( 20 ), internal_2_0( 20 ), internal_2_1( 21 ));
HA_16 : HA port map(internal_1_6( 20 ), internal_1_7( 20 ), internal_2_2( 20 ), internal_2_3( 21 ));
FA_44 : FA port map(internal_1_0( 21 ), internal_1_1( 21 ), internal_1_2( 21 ), internal_2_0( 21 ), internal_2_1( 22 ));
FA_45 : FA port map(internal_1_3( 21 ), internal_1_4( 21 ), internal_1_5( 21 ), internal_2_0( 21 ), internal_2_1( 22 ));
HA_17 : HA port map(internal_1_6( 21 ), internal_1_7( 21 ), internal_2_2( 21 ), internal_2_3( 22 ));
FA_46 : FA port map(internal_1_0( 22 ), internal_1_1( 22 ), internal_1_2( 22 ), internal_2_0( 22 ), internal_2_1( 23 ));
FA_47 : FA port map(internal_1_3( 22 ), internal_1_4( 22 ), internal_1_5( 22 ), internal_2_0( 22 ), internal_2_1( 23 ));
FA_48 : FA port map(internal_1_6( 22 ), internal_1_7( 22 ), internal_1_8( 22 ), internal_2_0( 22 ), internal_2_1( 23 ));
HA_18 : HA port map(internal_1_9( 22 ), internal_1_10( 22 ), internal_2_3( 22 ), internal_2_4( 23 ));
FA_49 : FA port map(internal_1_0( 23 ), internal_1_1( 23 ), internal_1_2( 23 ), internal_2_0( 23 ), internal_2_1( 24 ));
FA_50 : FA port map(internal_1_3( 23 ), internal_1_4( 23 ), internal_1_5( 23 ), internal_2_0( 23 ), internal_2_1( 24 ));
FA_51 : FA port map(internal_1_6( 23 ), internal_1_7( 23 ), internal_1_8( 23 ), internal_2_0( 23 ), internal_2_1( 24 ));
HA_19 : HA port map(internal_1_9( 23 ), internal_1_10( 23 ), internal_2_3( 23 ), internal_2_4( 24 ));
FA_52 : FA port map(internal_1_0( 24 ), internal_1_1( 24 ), internal_1_2( 24 ), internal_2_0( 24 ), internal_2_1( 25 ));
FA_53 : FA port map(internal_1_3( 24 ), internal_1_4( 24 ), internal_1_5( 24 ), internal_2_0( 24 ), internal_2_1( 25 ));
FA_54 : FA port map(internal_1_6( 24 ), internal_1_7( 24 ), internal_1_8( 24 ), internal_2_0( 24 ), internal_2_1( 25 ));
FA_55 : FA port map(internal_1_9( 24 ), internal_1_10( 24 ), internal_1_11( 24 ), internal_2_1( 24 ), internal_2_2( 25 ));
FA_56 : FA port map(internal_1_0( 25 ), internal_1_1( 25 ), internal_1_2( 25 ), internal_2_0( 25 ), internal_2_1( 26 ));
FA_57 : FA port map(internal_1_3( 25 ), internal_1_4( 25 ), internal_1_5( 25 ), internal_2_0( 25 ), internal_2_1( 26 ));
FA_58 : FA port map(internal_1_6( 25 ), internal_1_7( 25 ), internal_1_8( 25 ), internal_2_0( 25 ), internal_2_1( 26 ));
FA_59 : FA port map(internal_1_9( 25 ), internal_1_10( 25 ), internal_1_11( 25 ), internal_2_1( 25 ), internal_2_2( 26 ));
FA_60 : FA port map(internal_1_0( 26 ), internal_1_1( 26 ), internal_1_2( 26 ), internal_2_0( 26 ), internal_2_1( 27 ));
FA_61 : FA port map(internal_1_3( 26 ), internal_1_4( 26 ), internal_1_5( 26 ), internal_2_0( 26 ), internal_2_1( 27 ));
FA_62 : FA port map(internal_1_6( 26 ), internal_1_7( 26 ), internal_1_8( 26 ), internal_2_0( 26 ), internal_2_1( 27 ));
FA_63 : FA port map(internal_1_9( 26 ), internal_1_10( 26 ), internal_1_11( 26 ), internal_2_1( 26 ), internal_2_2( 27 ));
FA_64 : FA port map(internal_1_0( 27 ), internal_1_1( 27 ), internal_1_2( 27 ), internal_2_0( 27 ), internal_2_1( 28 ));
FA_65 : FA port map(internal_1_3( 27 ), internal_1_4( 27 ), internal_1_5( 27 ), internal_2_0( 27 ), internal_2_1( 28 ));
FA_66 : FA port map(internal_1_6( 27 ), internal_1_7( 27 ), internal_1_8( 27 ), internal_2_0( 27 ), internal_2_1( 28 ));
FA_67 : FA port map(internal_1_9( 27 ), internal_1_10( 27 ), internal_1_11( 27 ), internal_2_1( 27 ), internal_2_2( 28 ));
FA_68 : FA port map(internal_1_0( 28 ), internal_1_1( 28 ), internal_1_2( 28 ), internal_2_0( 28 ), internal_2_1( 29 ));
FA_69 : FA port map(internal_1_3( 28 ), internal_1_4( 28 ), internal_1_5( 28 ), internal_2_0( 28 ), internal_2_1( 29 ));
FA_70 : FA port map(internal_1_6( 28 ), internal_1_7( 28 ), internal_1_8( 28 ), internal_2_0( 28 ), internal_2_1( 29 ));
FA_71 : FA port map(internal_1_9( 28 ), internal_1_10( 28 ), internal_1_11( 28 ), internal_2_1( 28 ), internal_2_2( 29 ));
FA_72 : FA port map(internal_1_0( 29 ), internal_1_1( 29 ), internal_1_2( 29 ), internal_2_0( 29 ), internal_2_1( 30 ));
FA_73 : FA port map(internal_1_3( 29 ), internal_1_4( 29 ), internal_1_5( 29 ), internal_2_0( 29 ), internal_2_1( 30 ));
FA_74 : FA port map(internal_1_6( 29 ), internal_1_7( 29 ), internal_1_8( 29 ), internal_2_0( 29 ), internal_2_1( 30 ));
FA_75 : FA port map(internal_1_9( 29 ), internal_1_10( 29 ), internal_1_11( 29 ), internal_2_1( 29 ), internal_2_2( 30 ));
FA_76 : FA port map(internal_1_0( 30 ), internal_1_1( 30 ), internal_1_2( 30 ), internal_2_0( 30 ), internal_2_1( 31 ));
FA_77 : FA port map(internal_1_3( 30 ), internal_1_4( 30 ), internal_1_5( 30 ), internal_2_0( 30 ), internal_2_1( 31 ));
FA_78 : FA port map(internal_1_6( 30 ), internal_1_7( 30 ), internal_1_8( 30 ), internal_2_0( 30 ), internal_2_1( 31 ));
FA_79 : FA port map(internal_1_9( 30 ), internal_1_10( 30 ), internal_1_11( 30 ), internal_2_1( 30 ), internal_2_2( 31 ));
FA_80 : FA port map(internal_1_0( 31 ), internal_1_1( 31 ), internal_1_2( 31 ), internal_2_0( 31 ), internal_2_1( 32 ));
FA_81 : FA port map(internal_1_3( 31 ), internal_1_4( 31 ), internal_1_5( 31 ), internal_2_0( 31 ), internal_2_1( 32 ));
FA_82 : FA port map(internal_1_6( 31 ), internal_1_7( 31 ), internal_1_8( 31 ), internal_2_0( 31 ), internal_2_1( 32 ));
FA_83 : FA port map(internal_1_9( 31 ), internal_1_10( 31 ), internal_1_11( 31 ), internal_2_1( 31 ), internal_2_2( 32 ));
FA_84 : FA port map(internal_1_0( 32 ), internal_1_1( 32 ), internal_1_2( 32 ), internal_2_0( 32 ), internal_2_1( 33 ));
FA_85 : FA port map(internal_1_3( 32 ), internal_1_4( 32 ), internal_1_5( 32 ), internal_2_0( 32 ), internal_2_1( 33 ));
FA_86 : FA port map(internal_1_6( 32 ), internal_1_7( 32 ), internal_1_8( 32 ), internal_2_0( 32 ), internal_2_1( 33 ));
FA_87 : FA port map(internal_1_9( 32 ), internal_1_10( 32 ), internal_1_11( 32 ), internal_2_1( 32 ), internal_2_2( 33 ));
FA_88 : FA port map(internal_1_0( 33 ), internal_1_1( 33 ), internal_1_2( 33 ), internal_2_0( 33 ), internal_2_1( 34 ));
FA_89 : FA port map(internal_1_3( 33 ), internal_1_4( 33 ), internal_1_5( 33 ), internal_2_0( 33 ), internal_2_1( 34 ));
FA_90 : FA port map(internal_1_6( 33 ), internal_1_7( 33 ), internal_1_8( 33 ), internal_2_0( 33 ), internal_2_1( 34 ));
FA_91 : FA port map(internal_1_9( 33 ), internal_1_10( 33 ), internal_1_11( 33 ), internal_2_1( 33 ), internal_2_2( 34 ));
FA_92 : FA port map(internal_1_0( 34 ), internal_1_1( 34 ), internal_1_2( 34 ), internal_2_0( 34 ), internal_2_1( 35 ));
FA_93 : FA port map(internal_1_3( 34 ), internal_1_4( 34 ), internal_1_5( 34 ), internal_2_0( 34 ), internal_2_1( 35 ));
FA_94 : FA port map(internal_1_6( 34 ), internal_1_7( 34 ), internal_1_8( 34 ), internal_2_0( 34 ), internal_2_1( 35 ));
FA_95 : FA port map(internal_1_9( 34 ), internal_1_10( 34 ), internal_1_11( 34 ), internal_2_1( 34 ), internal_2_2( 35 ));
FA_96 : FA port map(internal_1_0( 35 ), internal_1_1( 35 ), internal_1_2( 35 ), internal_2_0( 35 ), internal_2_1( 36 ));
FA_97 : FA port map(internal_1_3( 35 ), internal_1_4( 35 ), internal_1_5( 35 ), internal_2_0( 35 ), internal_2_1( 36 ));
FA_98 : FA port map(internal_1_6( 35 ), internal_1_7( 35 ), internal_1_8( 35 ), internal_2_0( 35 ), internal_2_1( 36 ));
FA_99 : FA port map(internal_1_9( 35 ), internal_1_10( 35 ), internal_1_11( 35 ), internal_2_1( 35 ), internal_2_2( 36 ));
FA_100 : FA port map(internal_1_0( 36 ), internal_1_1( 36 ), internal_1_2( 36 ), internal_2_0( 36 ), internal_2_1( 37 ));
FA_101 : FA port map(internal_1_3( 36 ), internal_1_4( 36 ), internal_1_5( 36 ), internal_2_0( 36 ), internal_2_1( 37 ));
FA_102 : FA port map(internal_1_6( 36 ), internal_1_7( 36 ), internal_1_8( 36 ), internal_2_0( 36 ), internal_2_1( 37 ));
FA_103 : FA port map(internal_1_9( 36 ), internal_1_10( 36 ), internal_1_11( 36 ), internal_2_1( 36 ), internal_2_2( 37 ));
FA_104 : FA port map(internal_1_0( 37 ), internal_1_1( 37 ), internal_1_2( 37 ), internal_2_0( 37 ), internal_2_1( 38 ));
FA_105 : FA port map(internal_1_3( 37 ), internal_1_4( 37 ), internal_1_5( 37 ), internal_2_0( 37 ), internal_2_1( 38 ));
FA_106 : FA port map(internal_1_6( 37 ), internal_1_7( 37 ), internal_1_8( 37 ), internal_2_0( 37 ), internal_2_1( 38 ));
FA_107 : FA port map(internal_1_9( 37 ), internal_1_10( 37 ), internal_1_11( 37 ), internal_2_1( 37 ), internal_2_2( 38 ));
FA_108 : FA port map(internal_1_0( 38 ), internal_1_1( 38 ), internal_1_2( 38 ), internal_2_0( 38 ), internal_2_1( 39 ));
FA_109 : FA port map(internal_1_3( 38 ), internal_1_4( 38 ), internal_1_5( 38 ), internal_2_0( 38 ), internal_2_1( 39 ));
FA_110 : FA port map(internal_1_6( 38 ), internal_1_7( 38 ), internal_1_8( 38 ), internal_2_0( 38 ), internal_2_1( 39 ));
FA_111 : FA port map(internal_1_9( 38 ), internal_1_10( 38 ), internal_1_11( 38 ), internal_2_1( 38 ), internal_2_2( 39 ));
FA_112 : FA port map(internal_1_0( 39 ), internal_1_1( 39 ), internal_1_2( 39 ), internal_2_0( 39 ), internal_2_1( 40 ));
FA_113 : FA port map(internal_1_3( 39 ), internal_1_4( 39 ), internal_1_5( 39 ), internal_2_0( 39 ), internal_2_1( 40 ));
FA_114 : FA port map(internal_1_6( 39 ), internal_1_7( 39 ), internal_1_8( 39 ), internal_2_0( 39 ), internal_2_1( 40 ));
FA_115 : FA port map(internal_1_9( 39 ), internal_1_10( 39 ), internal_1_11( 39 ), internal_2_1( 39 ), internal_2_2( 40 ));
FA_116 : FA port map(internal_1_0( 40 ), internal_1_1( 40 ), internal_1_2( 40 ), internal_2_0( 40 ), internal_2_1( 41 ));
FA_117 : FA port map(internal_1_3( 40 ), internal_1_4( 40 ), internal_1_5( 40 ), internal_2_0( 40 ), internal_2_1( 41 ));
FA_118 : FA port map(internal_1_6( 40 ), internal_1_7( 40 ), internal_1_8( 40 ), internal_2_0( 40 ), internal_2_1( 41 ));
FA_119 : FA port map(internal_1_9( 40 ), internal_1_10( 40 ), internal_1_11( 40 ), internal_2_1( 40 ), internal_2_2( 41 ));
FA_120 : FA port map(internal_1_0( 41 ), internal_1_1( 41 ), internal_1_2( 41 ), internal_2_0( 41 ), internal_2_1( 42 ));
FA_121 : FA port map(internal_1_3( 41 ), internal_1_4( 41 ), internal_1_5( 41 ), internal_2_0( 41 ), internal_2_1( 42 ));
FA_122 : FA port map(internal_1_6( 41 ), internal_1_7( 41 ), internal_1_8( 41 ), internal_2_0( 41 ), internal_2_1( 42 ));
FA_123 : FA port map(internal_1_9( 41 ), internal_1_10( 41 ), internal_1_11( 41 ), internal_2_1( 41 ), internal_2_2( 42 ));
FA_124 : FA port map(internal_1_0( 42 ), internal_1_1( 42 ), internal_1_2( 42 ), internal_2_0( 42 ), internal_2_1( 43 ));
FA_125 : FA port map(internal_1_3( 42 ), internal_1_4( 42 ), internal_1_5( 42 ), internal_2_0( 42 ), internal_2_1( 43 ));
FA_126 : FA port map(internal_1_6( 42 ), internal_1_7( 42 ), internal_1_8( 42 ), internal_2_0( 42 ), internal_2_1( 43 ));
FA_127 : FA port map(internal_1_9( 42 ), internal_1_10( 42 ), internal_1_11( 42 ), internal_2_1( 42 ), internal_2_2( 43 ));
FA_128 : FA port map(internal_1_0( 43 ), internal_1_1( 43 ), internal_1_2( 43 ), internal_2_0( 43 ), internal_2_1( 44 ));
FA_129 : FA port map(internal_1_3( 43 ), internal_1_4( 43 ), internal_1_5( 43 ), internal_2_0( 43 ), internal_2_1( 44 ));
FA_130 : FA port map(internal_1_6( 43 ), internal_1_7( 43 ), internal_1_8( 43 ), internal_2_0( 43 ), internal_2_1( 44 ));
HA_20 : HA port map(internal_1_9( 43 ), internal_1_10( 43 ), internal_2_3( 43 ), internal_2_4( 44 ));
FA_131 : FA port map(internal_1_0( 44 ), internal_1_1( 44 ), internal_1_2( 44 ), internal_2_0( 44 ), internal_2_1( 45 ));
FA_132 : FA port map(internal_1_3( 44 ), internal_1_4( 44 ), internal_1_5( 44 ), internal_2_0( 44 ), internal_2_1( 45 ));
FA_133 : FA port map(internal_1_6( 44 ), internal_1_7( 44 ), internal_1_8( 44 ), internal_2_0( 44 ), internal_2_1( 45 ));
HA_21 : HA port map(internal_1_9( 44 ), internal_1_10( 44 ), internal_2_3( 44 ), internal_2_4( 45 ));
FA_134 : FA port map(internal_1_0( 45 ), internal_1_1( 45 ), internal_1_2( 45 ), internal_2_0( 45 ), internal_2_1( 46 ));
FA_135 : FA port map(internal_1_3( 45 ), internal_1_4( 45 ), internal_1_5( 45 ), internal_2_0( 45 ), internal_2_1( 46 ));
FA_136 : FA port map(internal_1_6( 45 ), internal_1_7( 45 ), internal_1_8( 45 ), internal_2_0( 45 ), internal_2_1( 46 ));
FA_137 : FA port map(internal_1_0( 46 ), internal_1_1( 46 ), internal_1_2( 46 ), internal_2_0( 46 ), internal_2_1( 47 ));
FA_138 : FA port map(internal_1_3( 46 ), internal_1_4( 46 ), internal_1_5( 46 ), internal_2_0( 46 ), internal_2_1( 47 ));
HA_22 : HA port map(internal_1_6( 46 ), internal_1_7( 46 ), internal_2_2( 46 ), internal_2_3( 47 ));
FA_139 : FA port map(internal_1_0( 47 ), internal_1_1( 47 ), internal_1_2( 47 ), internal_2_0( 47 ), internal_2_1( 48 ));
FA_140 : FA port map(internal_1_3( 47 ), internal_1_4( 47 ), internal_1_5( 47 ), internal_2_0( 47 ), internal_2_1( 48 ));
FA_141 : FA port map(internal_1_0( 48 ), internal_1_1( 48 ), internal_1_2( 48 ), internal_2_0( 48 ), internal_2_1( 49 ));
HA_23 : HA port map(internal_1_3( 48 ), internal_1_4( 48 ), internal_2_1( 48 ), internal_2_2( 49 ));
FA_142 : FA port map(internal_1_0( 49 ), internal_1_1( 49 ), internal_1_2( 49 ), internal_2_0( 49 ), internal_2_1( 50 ));
HA_24 : HA port map(internal_1_0( 50 ), internal_1_1( 50 ), internal_2_0( 50 ), internal_2_1( 51 ));
HA_25 : HA port map(internal_2_0( 10 ), internal_2_1( 10 ), internal_3_0( 10 ), internal_3_1( 11 ));
HA_26 : HA port map(internal_2_0( 11 ), internal_2_1( 11 ), internal_3_0( 11 ), internal_3_1( 12 ));
FA_143 : FA port map(internal_2_0( 12 ), internal_2_1( 12 ), internal_2_2( 12 ), internal_3_0( 12 ), internal_3_1( 13 ));
HA_27 : HA port map(internal_2_3( 12 ), internal_2_4( 12 ), internal_3_1( 12 ), internal_3_2( 13 ));
FA_144 : FA port map(internal_2_0( 13 ), internal_2_1( 13 ), internal_2_2( 13 ), internal_3_0( 13 ), internal_3_1( 14 ));
HA_28 : HA port map(internal_2_3( 13 ), internal_2_4( 13 ), internal_3_1( 13 ), internal_3_2( 14 ));
FA_145 : FA port map(internal_2_0( 14 ), internal_2_1( 14 ), internal_2_2( 14 ), internal_3_0( 14 ), internal_3_1( 15 ));
FA_146 : FA port map(internal_2_3( 14 ), internal_2_4( 14 ), internal_2_5( 14 ), internal_3_0( 14 ), internal_3_1( 15 ));
HA_29 : HA port map(internal_2_6( 14 ), internal_2_7( 14 ), internal_3_2( 14 ), internal_3_3( 15 ));
FA_147 : FA port map(internal_2_0( 15 ), internal_2_1( 15 ), internal_2_2( 15 ), internal_3_0( 15 ), internal_3_1( 16 ));
FA_148 : FA port map(internal_2_3( 15 ), internal_2_4( 15 ), internal_2_5( 15 ), internal_3_0( 15 ), internal_3_1( 16 ));
HA_30 : HA port map(internal_2_6( 15 ), internal_2_7( 15 ), internal_3_2( 15 ), internal_3_3( 16 ));
FA_149 : FA port map(internal_2_0( 16 ), internal_2_1( 16 ), internal_2_2( 16 ), internal_3_0( 16 ), internal_3_1( 17 ));
FA_150 : FA port map(internal_2_3( 16 ), internal_2_4( 16 ), internal_2_5( 16 ), internal_3_0( 16 ), internal_3_1( 17 ));
FA_151 : FA port map(internal_2_6( 16 ), internal_2_7( 16 ), internal_2_8( 16 ), internal_3_0( 16 ), internal_3_1( 17 ));
FA_152 : FA port map(internal_2_0( 17 ), internal_2_1( 17 ), internal_2_2( 17 ), internal_3_0( 17 ), internal_3_1( 18 ));
FA_153 : FA port map(internal_2_3( 17 ), internal_2_4( 17 ), internal_2_5( 17 ), internal_3_0( 17 ), internal_3_1( 18 ));
FA_154 : FA port map(internal_2_6( 17 ), internal_2_7( 17 ), internal_2_8( 17 ), internal_3_0( 17 ), internal_3_1( 18 ));
FA_155 : FA port map(internal_2_0( 18 ), internal_2_1( 18 ), internal_2_2( 18 ), internal_3_0( 18 ), internal_3_1( 19 ));
FA_156 : FA port map(internal_2_3( 18 ), internal_2_4( 18 ), internal_2_5( 18 ), internal_3_0( 18 ), internal_3_1( 19 ));
FA_157 : FA port map(internal_2_6( 18 ), internal_2_7( 18 ), internal_2_8( 18 ), internal_3_0( 18 ), internal_3_1( 19 ));
FA_158 : FA port map(internal_2_0( 19 ), internal_2_1( 19 ), internal_2_2( 19 ), internal_3_0( 19 ), internal_3_1( 20 ));
FA_159 : FA port map(internal_2_3( 19 ), internal_2_4( 19 ), internal_2_5( 19 ), internal_3_0( 19 ), internal_3_1( 20 ));
FA_160 : FA port map(internal_2_6( 19 ), internal_2_7( 19 ), internal_2_8( 19 ), internal_3_0( 19 ), internal_3_1( 20 ));
FA_161 : FA port map(internal_2_0( 20 ), internal_2_1( 20 ), internal_2_2( 20 ), internal_3_0( 20 ), internal_3_1( 21 ));
FA_162 : FA port map(internal_2_3( 20 ), internal_2_4( 20 ), internal_2_5( 20 ), internal_3_0( 20 ), internal_3_1( 21 ));
FA_163 : FA port map(internal_2_6( 20 ), internal_2_7( 20 ), internal_2_8( 20 ), internal_3_0( 20 ), internal_3_1( 21 ));
FA_164 : FA port map(internal_2_0( 21 ), internal_2_1( 21 ), internal_2_2( 21 ), internal_3_0( 21 ), internal_3_1( 22 ));
FA_165 : FA port map(internal_2_3( 21 ), internal_2_4( 21 ), internal_2_5( 21 ), internal_3_0( 21 ), internal_3_1( 22 ));
FA_166 : FA port map(internal_2_6( 21 ), internal_2_7( 21 ), internal_2_8( 21 ), internal_3_0( 21 ), internal_3_1( 22 ));
FA_167 : FA port map(internal_2_0( 22 ), internal_2_1( 22 ), internal_2_2( 22 ), internal_3_0( 22 ), internal_3_1( 23 ));
FA_168 : FA port map(internal_2_3( 22 ), internal_2_4( 22 ), internal_2_5( 22 ), internal_3_0( 22 ), internal_3_1( 23 ));
FA_169 : FA port map(internal_2_6( 22 ), internal_2_7( 22 ), internal_2_8( 22 ), internal_3_0( 22 ), internal_3_1( 23 ));
FA_170 : FA port map(internal_2_0( 23 ), internal_2_1( 23 ), internal_2_2( 23 ), internal_3_0( 23 ), internal_3_1( 24 ));
FA_171 : FA port map(internal_2_3( 23 ), internal_2_4( 23 ), internal_2_5( 23 ), internal_3_0( 23 ), internal_3_1( 24 ));
FA_172 : FA port map(internal_2_6( 23 ), internal_2_7( 23 ), internal_2_8( 23 ), internal_3_0( 23 ), internal_3_1( 24 ));
FA_173 : FA port map(internal_2_0( 24 ), internal_2_1( 24 ), internal_2_2( 24 ), internal_3_0( 24 ), internal_3_1( 25 ));
FA_174 : FA port map(internal_2_3( 24 ), internal_2_4( 24 ), internal_2_5( 24 ), internal_3_0( 24 ), internal_3_1( 25 ));
FA_175 : FA port map(internal_2_6( 24 ), internal_2_7( 24 ), internal_2_8( 24 ), internal_3_0( 24 ), internal_3_1( 25 ));
FA_176 : FA port map(internal_2_0( 25 ), internal_2_1( 25 ), internal_2_2( 25 ), internal_3_0( 25 ), internal_3_1( 26 ));
FA_177 : FA port map(internal_2_3( 25 ), internal_2_4( 25 ), internal_2_5( 25 ), internal_3_0( 25 ), internal_3_1( 26 ));
FA_178 : FA port map(internal_2_6( 25 ), internal_2_7( 25 ), internal_2_8( 25 ), internal_3_0( 25 ), internal_3_1( 26 ));
FA_179 : FA port map(internal_2_0( 26 ), internal_2_1( 26 ), internal_2_2( 26 ), internal_3_0( 26 ), internal_3_1( 27 ));
FA_180 : FA port map(internal_2_3( 26 ), internal_2_4( 26 ), internal_2_5( 26 ), internal_3_0( 26 ), internal_3_1( 27 ));
FA_181 : FA port map(internal_2_6( 26 ), internal_2_7( 26 ), internal_2_8( 26 ), internal_3_0( 26 ), internal_3_1( 27 ));
FA_182 : FA port map(internal_2_0( 27 ), internal_2_1( 27 ), internal_2_2( 27 ), internal_3_0( 27 ), internal_3_1( 28 ));
FA_183 : FA port map(internal_2_3( 27 ), internal_2_4( 27 ), internal_2_5( 27 ), internal_3_0( 27 ), internal_3_1( 28 ));
FA_184 : FA port map(internal_2_6( 27 ), internal_2_7( 27 ), internal_2_8( 27 ), internal_3_0( 27 ), internal_3_1( 28 ));
FA_185 : FA port map(internal_2_0( 28 ), internal_2_1( 28 ), internal_2_2( 28 ), internal_3_0( 28 ), internal_3_1( 29 ));
FA_186 : FA port map(internal_2_3( 28 ), internal_2_4( 28 ), internal_2_5( 28 ), internal_3_0( 28 ), internal_3_1( 29 ));
FA_187 : FA port map(internal_2_6( 28 ), internal_2_7( 28 ), internal_2_8( 28 ), internal_3_0( 28 ), internal_3_1( 29 ));
FA_188 : FA port map(internal_2_0( 29 ), internal_2_1( 29 ), internal_2_2( 29 ), internal_3_0( 29 ), internal_3_1( 30 ));
FA_189 : FA port map(internal_2_3( 29 ), internal_2_4( 29 ), internal_2_5( 29 ), internal_3_0( 29 ), internal_3_1( 30 ));
FA_190 : FA port map(internal_2_6( 29 ), internal_2_7( 29 ), internal_2_8( 29 ), internal_3_0( 29 ), internal_3_1( 30 ));
FA_191 : FA port map(internal_2_0( 30 ), internal_2_1( 30 ), internal_2_2( 30 ), internal_3_0( 30 ), internal_3_1( 31 ));
FA_192 : FA port map(internal_2_3( 30 ), internal_2_4( 30 ), internal_2_5( 30 ), internal_3_0( 30 ), internal_3_1( 31 ));
FA_193 : FA port map(internal_2_6( 30 ), internal_2_7( 30 ), internal_2_8( 30 ), internal_3_0( 30 ), internal_3_1( 31 ));
FA_194 : FA port map(internal_2_0( 31 ), internal_2_1( 31 ), internal_2_2( 31 ), internal_3_0( 31 ), internal_3_1( 32 ));
FA_195 : FA port map(internal_2_3( 31 ), internal_2_4( 31 ), internal_2_5( 31 ), internal_3_0( 31 ), internal_3_1( 32 ));
FA_196 : FA port map(internal_2_6( 31 ), internal_2_7( 31 ), internal_2_8( 31 ), internal_3_0( 31 ), internal_3_1( 32 ));
FA_197 : FA port map(internal_2_0( 32 ), internal_2_1( 32 ), internal_2_2( 32 ), internal_3_0( 32 ), internal_3_1( 33 ));
FA_198 : FA port map(internal_2_3( 32 ), internal_2_4( 32 ), internal_2_5( 32 ), internal_3_0( 32 ), internal_3_1( 33 ));
FA_199 : FA port map(internal_2_6( 32 ), internal_2_7( 32 ), internal_2_8( 32 ), internal_3_0( 32 ), internal_3_1( 33 ));
FA_200 : FA port map(internal_2_0( 33 ), internal_2_1( 33 ), internal_2_2( 33 ), internal_3_0( 33 ), internal_3_1( 34 ));
FA_201 : FA port map(internal_2_3( 33 ), internal_2_4( 33 ), internal_2_5( 33 ), internal_3_0( 33 ), internal_3_1( 34 ));
FA_202 : FA port map(internal_2_6( 33 ), internal_2_7( 33 ), internal_2_8( 33 ), internal_3_0( 33 ), internal_3_1( 34 ));
FA_203 : FA port map(internal_2_0( 34 ), internal_2_1( 34 ), internal_2_2( 34 ), internal_3_0( 34 ), internal_3_1( 35 ));
FA_204 : FA port map(internal_2_3( 34 ), internal_2_4( 34 ), internal_2_5( 34 ), internal_3_0( 34 ), internal_3_1( 35 ));
FA_205 : FA port map(internal_2_6( 34 ), internal_2_7( 34 ), internal_2_8( 34 ), internal_3_0( 34 ), internal_3_1( 35 ));
FA_206 : FA port map(internal_2_0( 35 ), internal_2_1( 35 ), internal_2_2( 35 ), internal_3_0( 35 ), internal_3_1( 36 ));
FA_207 : FA port map(internal_2_3( 35 ), internal_2_4( 35 ), internal_2_5( 35 ), internal_3_0( 35 ), internal_3_1( 36 ));
FA_208 : FA port map(internal_2_6( 35 ), internal_2_7( 35 ), internal_2_8( 35 ), internal_3_0( 35 ), internal_3_1( 36 ));
FA_209 : FA port map(internal_2_0( 36 ), internal_2_1( 36 ), internal_2_2( 36 ), internal_3_0( 36 ), internal_3_1( 37 ));
FA_210 : FA port map(internal_2_3( 36 ), internal_2_4( 36 ), internal_2_5( 36 ), internal_3_0( 36 ), internal_3_1( 37 ));
FA_211 : FA port map(internal_2_6( 36 ), internal_2_7( 36 ), internal_2_8( 36 ), internal_3_0( 36 ), internal_3_1( 37 ));
FA_212 : FA port map(internal_2_0( 37 ), internal_2_1( 37 ), internal_2_2( 37 ), internal_3_0( 37 ), internal_3_1( 38 ));
FA_213 : FA port map(internal_2_3( 37 ), internal_2_4( 37 ), internal_2_5( 37 ), internal_3_0( 37 ), internal_3_1( 38 ));
FA_214 : FA port map(internal_2_6( 37 ), internal_2_7( 37 ), internal_2_8( 37 ), internal_3_0( 37 ), internal_3_1( 38 ));
FA_215 : FA port map(internal_2_0( 38 ), internal_2_1( 38 ), internal_2_2( 38 ), internal_3_0( 38 ), internal_3_1( 39 ));
FA_216 : FA port map(internal_2_3( 38 ), internal_2_4( 38 ), internal_2_5( 38 ), internal_3_0( 38 ), internal_3_1( 39 ));
FA_217 : FA port map(internal_2_6( 38 ), internal_2_7( 38 ), internal_2_8( 38 ), internal_3_0( 38 ), internal_3_1( 39 ));
FA_218 : FA port map(internal_2_0( 39 ), internal_2_1( 39 ), internal_2_2( 39 ), internal_3_0( 39 ), internal_3_1( 40 ));
FA_219 : FA port map(internal_2_3( 39 ), internal_2_4( 39 ), internal_2_5( 39 ), internal_3_0( 39 ), internal_3_1( 40 ));
FA_220 : FA port map(internal_2_6( 39 ), internal_2_7( 39 ), internal_2_8( 39 ), internal_3_0( 39 ), internal_3_1( 40 ));
FA_221 : FA port map(internal_2_0( 40 ), internal_2_1( 40 ), internal_2_2( 40 ), internal_3_0( 40 ), internal_3_1( 41 ));
FA_222 : FA port map(internal_2_3( 40 ), internal_2_4( 40 ), internal_2_5( 40 ), internal_3_0( 40 ), internal_3_1( 41 ));
FA_223 : FA port map(internal_2_6( 40 ), internal_2_7( 40 ), internal_2_8( 40 ), internal_3_0( 40 ), internal_3_1( 41 ));
FA_224 : FA port map(internal_2_0( 41 ), internal_2_1( 41 ), internal_2_2( 41 ), internal_3_0( 41 ), internal_3_1( 42 ));
FA_225 : FA port map(internal_2_3( 41 ), internal_2_4( 41 ), internal_2_5( 41 ), internal_3_0( 41 ), internal_3_1( 42 ));
FA_226 : FA port map(internal_2_6( 41 ), internal_2_7( 41 ), internal_2_8( 41 ), internal_3_0( 41 ), internal_3_1( 42 ));
FA_227 : FA port map(internal_2_0( 42 ), internal_2_1( 42 ), internal_2_2( 42 ), internal_3_0( 42 ), internal_3_1( 43 ));
FA_228 : FA port map(internal_2_3( 42 ), internal_2_4( 42 ), internal_2_5( 42 ), internal_3_0( 42 ), internal_3_1( 43 ));
FA_229 : FA port map(internal_2_6( 42 ), internal_2_7( 42 ), internal_2_8( 42 ), internal_3_0( 42 ), internal_3_1( 43 ));
FA_230 : FA port map(internal_2_0( 43 ), internal_2_1( 43 ), internal_2_2( 43 ), internal_3_0( 43 ), internal_3_1( 44 ));
FA_231 : FA port map(internal_2_3( 43 ), internal_2_4( 43 ), internal_2_5( 43 ), internal_3_0( 43 ), internal_3_1( 44 ));
FA_232 : FA port map(internal_2_6( 43 ), internal_2_7( 43 ), internal_2_8( 43 ), internal_3_0( 43 ), internal_3_1( 44 ));
FA_233 : FA port map(internal_2_0( 44 ), internal_2_1( 44 ), internal_2_2( 44 ), internal_3_0( 44 ), internal_3_1( 45 ));
FA_234 : FA port map(internal_2_3( 44 ), internal_2_4( 44 ), internal_2_5( 44 ), internal_3_0( 44 ), internal_3_1( 45 ));
FA_235 : FA port map(internal_2_6( 44 ), internal_2_7( 44 ), internal_2_8( 44 ), internal_3_0( 44 ), internal_3_1( 45 ));
FA_236 : FA port map(internal_2_0( 45 ), internal_2_1( 45 ), internal_2_2( 45 ), internal_3_0( 45 ), internal_3_1( 46 ));
FA_237 : FA port map(internal_2_3( 45 ), internal_2_4( 45 ), internal_2_5( 45 ), internal_3_0( 45 ), internal_3_1( 46 ));
FA_238 : FA port map(internal_2_6( 45 ), internal_2_7( 45 ), internal_2_8( 45 ), internal_3_0( 45 ), internal_3_1( 46 ));
FA_239 : FA port map(internal_2_0( 46 ), internal_2_1( 46 ), internal_2_2( 46 ), internal_3_0( 46 ), internal_3_1( 47 ));
FA_240 : FA port map(internal_2_3( 46 ), internal_2_4( 46 ), internal_2_5( 46 ), internal_3_0( 46 ), internal_3_1( 47 ));
FA_241 : FA port map(internal_2_6( 46 ), internal_2_7( 46 ), internal_2_8( 46 ), internal_3_0( 46 ), internal_3_1( 47 ));
FA_242 : FA port map(internal_2_0( 47 ), internal_2_1( 47 ), internal_2_2( 47 ), internal_3_0( 47 ), internal_3_1( 48 ));
FA_243 : FA port map(internal_2_3( 47 ), internal_2_4( 47 ), internal_2_5( 47 ), internal_3_0( 47 ), internal_3_1( 48 ));
FA_244 : FA port map(internal_2_6( 47 ), internal_2_7( 47 ), internal_2_8( 47 ), internal_3_0( 47 ), internal_3_1( 48 ));
FA_245 : FA port map(internal_2_0( 48 ), internal_2_1( 48 ), internal_2_2( 48 ), internal_3_0( 48 ), internal_3_1( 49 ));
FA_246 : FA port map(internal_2_3( 48 ), internal_2_4( 48 ), internal_2_5( 48 ), internal_3_0( 48 ), internal_3_1( 49 ));
FA_247 : FA port map(internal_2_6( 48 ), internal_2_7( 48 ), internal_2_8( 48 ), internal_3_0( 48 ), internal_3_1( 49 ));
FA_248 : FA port map(internal_2_0( 49 ), internal_2_1( 49 ), internal_2_2( 49 ), internal_3_0( 49 ), internal_3_1( 50 ));
FA_249 : FA port map(internal_2_3( 49 ), internal_2_4( 49 ), internal_2_5( 49 ), internal_3_0( 49 ), internal_3_1( 50 ));
FA_250 : FA port map(internal_2_6( 49 ), internal_2_7( 49 ), internal_2_8( 49 ), internal_3_0( 49 ), internal_3_1( 50 ));
FA_251 : FA port map(internal_2_0( 50 ), internal_2_1( 50 ), internal_2_2( 50 ), internal_3_0( 50 ), internal_3_1( 51 ));
FA_252 : FA port map(internal_2_3( 50 ), internal_2_4( 50 ), internal_2_5( 50 ), internal_3_0( 50 ), internal_3_1( 51 ));
FA_253 : FA port map(internal_2_6( 50 ), internal_2_7( 50 ), internal_2_8( 50 ), internal_3_0( 50 ), internal_3_1( 51 ));
FA_254 : FA port map(internal_2_0( 51 ), internal_2_1( 51 ), internal_2_2( 51 ), internal_3_0( 51 ), internal_3_1( 52 ));
FA_255 : FA port map(internal_2_3( 51 ), internal_2_4( 51 ), internal_2_5( 51 ), internal_3_0( 51 ), internal_3_1( 52 ));
HA_31 : HA port map(internal_2_6( 51 ), internal_2_7( 51 ), internal_3_2( 51 ), internal_3_3( 52 ));
FA_256 : FA port map(internal_2_0( 52 ), internal_2_1( 52 ), internal_2_2( 52 ), internal_3_0( 52 ), internal_3_1( 53 ));
FA_257 : FA port map(internal_2_3( 52 ), internal_2_4( 52 ), internal_2_5( 52 ), internal_3_0( 52 ), internal_3_1( 53 ));
HA_32 : HA port map(internal_2_6( 52 ), internal_2_7( 52 ), internal_3_2( 52 ), internal_3_3( 53 ));
FA_258 : FA port map(internal_2_0( 53 ), internal_2_1( 53 ), internal_2_2( 53 ), internal_3_0( 53 ), internal_3_1( 54 ));
FA_259 : FA port map(internal_2_3( 53 ), internal_2_4( 53 ), internal_2_5( 53 ), internal_3_0( 53 ), internal_3_1( 54 ));
FA_260 : FA port map(internal_2_0( 54 ), internal_2_1( 54 ), internal_2_2( 54 ), internal_3_0( 54 ), internal_3_1( 55 ));
HA_33 : HA port map(internal_2_3( 54 ), internal_2_4( 54 ), internal_3_1( 54 ), internal_3_2( 55 ));
FA_261 : FA port map(internal_2_0( 55 ), internal_2_1( 55 ), internal_2_2( 55 ), internal_3_0( 55 ), internal_3_1( 56 ));
HA_34 : HA port map(internal_2_0( 56 ), internal_2_1( 56 ), internal_3_0( 56 ), internal_3_1( 57 ));
HA_35 : HA port map(internal_3_0( 6 ), internal_3_1( 6 ), internal_4_0( 6 ), internal_4_1( 7 ));
HA_36 : HA port map(internal_3_0( 7 ), internal_3_1( 7 ), internal_4_0( 7 ), internal_4_1( 8 ));
FA_262 : FA port map(internal_3_0( 8 ), internal_3_1( 8 ), internal_3_2( 8 ), internal_4_0( 8 ), internal_4_1( 9 ));
HA_37 : HA port map(internal_3_3( 8 ), internal_3_4( 8 ), internal_4_1( 8 ), internal_4_2( 9 ));
FA_263 : FA port map(internal_3_0( 9 ), internal_3_1( 9 ), internal_3_2( 9 ), internal_4_0( 9 ), internal_4_1( 10 ));
HA_38 : HA port map(internal_3_3( 9 ), internal_3_4( 9 ), internal_4_1( 9 ), internal_4_2( 10 ));
FA_264 : FA port map(internal_3_0( 10 ), internal_3_1( 10 ), internal_3_2( 10 ), internal_4_0( 10 ), internal_4_1( 11 ));
FA_265 : FA port map(internal_3_3( 10 ), internal_3_4( 10 ), internal_3_5( 10 ), internal_4_0( 10 ), internal_4_1( 11 ));
FA_266 : FA port map(internal_3_0( 11 ), internal_3_1( 11 ), internal_3_2( 11 ), internal_4_0( 11 ), internal_4_1( 12 ));
FA_267 : FA port map(internal_3_3( 11 ), internal_3_4( 11 ), internal_3_5( 11 ), internal_4_0( 11 ), internal_4_1( 12 ));
FA_268 : FA port map(internal_3_0( 12 ), internal_3_1( 12 ), internal_3_2( 12 ), internal_4_0( 12 ), internal_4_1( 13 ));
FA_269 : FA port map(internal_3_3( 12 ), internal_3_4( 12 ), internal_3_5( 12 ), internal_4_0( 12 ), internal_4_1( 13 ));
FA_270 : FA port map(internal_3_0( 13 ), internal_3_1( 13 ), internal_3_2( 13 ), internal_4_0( 13 ), internal_4_1( 14 ));
FA_271 : FA port map(internal_3_3( 13 ), internal_3_4( 13 ), internal_3_5( 13 ), internal_4_0( 13 ), internal_4_1( 14 ));
FA_272 : FA port map(internal_3_0( 14 ), internal_3_1( 14 ), internal_3_2( 14 ), internal_4_0( 14 ), internal_4_1( 15 ));
FA_273 : FA port map(internal_3_3( 14 ), internal_3_4( 14 ), internal_3_5( 14 ), internal_4_0( 14 ), internal_4_1( 15 ));
FA_274 : FA port map(internal_3_0( 15 ), internal_3_1( 15 ), internal_3_2( 15 ), internal_4_0( 15 ), internal_4_1( 16 ));
FA_275 : FA port map(internal_3_3( 15 ), internal_3_4( 15 ), internal_3_5( 15 ), internal_4_0( 15 ), internal_4_1( 16 ));
FA_276 : FA port map(internal_3_0( 16 ), internal_3_1( 16 ), internal_3_2( 16 ), internal_4_0( 16 ), internal_4_1( 17 ));
FA_277 : FA port map(internal_3_3( 16 ), internal_3_4( 16 ), internal_3_5( 16 ), internal_4_0( 16 ), internal_4_1( 17 ));
FA_278 : FA port map(internal_3_0( 17 ), internal_3_1( 17 ), internal_3_2( 17 ), internal_4_0( 17 ), internal_4_1( 18 ));
FA_279 : FA port map(internal_3_3( 17 ), internal_3_4( 17 ), internal_3_5( 17 ), internal_4_0( 17 ), internal_4_1( 18 ));
FA_280 : FA port map(internal_3_0( 18 ), internal_3_1( 18 ), internal_3_2( 18 ), internal_4_0( 18 ), internal_4_1( 19 ));
FA_281 : FA port map(internal_3_3( 18 ), internal_3_4( 18 ), internal_3_5( 18 ), internal_4_0( 18 ), internal_4_1( 19 ));
FA_282 : FA port map(internal_3_0( 19 ), internal_3_1( 19 ), internal_3_2( 19 ), internal_4_0( 19 ), internal_4_1( 20 ));
FA_283 : FA port map(internal_3_3( 19 ), internal_3_4( 19 ), internal_3_5( 19 ), internal_4_0( 19 ), internal_4_1( 20 ));
FA_284 : FA port map(internal_3_0( 20 ), internal_3_1( 20 ), internal_3_2( 20 ), internal_4_0( 20 ), internal_4_1( 21 ));
FA_285 : FA port map(internal_3_3( 20 ), internal_3_4( 20 ), internal_3_5( 20 ), internal_4_0( 20 ), internal_4_1( 21 ));
FA_286 : FA port map(internal_3_0( 21 ), internal_3_1( 21 ), internal_3_2( 21 ), internal_4_0( 21 ), internal_4_1( 22 ));
FA_287 : FA port map(internal_3_3( 21 ), internal_3_4( 21 ), internal_3_5( 21 ), internal_4_0( 21 ), internal_4_1( 22 ));
FA_288 : FA port map(internal_3_0( 22 ), internal_3_1( 22 ), internal_3_2( 22 ), internal_4_0( 22 ), internal_4_1( 23 ));
FA_289 : FA port map(internal_3_3( 22 ), internal_3_4( 22 ), internal_3_5( 22 ), internal_4_0( 22 ), internal_4_1( 23 ));
FA_290 : FA port map(internal_3_0( 23 ), internal_3_1( 23 ), internal_3_2( 23 ), internal_4_0( 23 ), internal_4_1( 24 ));
FA_291 : FA port map(internal_3_3( 23 ), internal_3_4( 23 ), internal_3_5( 23 ), internal_4_0( 23 ), internal_4_1( 24 ));
FA_292 : FA port map(internal_3_0( 24 ), internal_3_1( 24 ), internal_3_2( 24 ), internal_4_0( 24 ), internal_4_1( 25 ));
FA_293 : FA port map(internal_3_3( 24 ), internal_3_4( 24 ), internal_3_5( 24 ), internal_4_0( 24 ), internal_4_1( 25 ));
FA_294 : FA port map(internal_3_0( 25 ), internal_3_1( 25 ), internal_3_2( 25 ), internal_4_0( 25 ), internal_4_1( 26 ));
FA_295 : FA port map(internal_3_3( 25 ), internal_3_4( 25 ), internal_3_5( 25 ), internal_4_0( 25 ), internal_4_1( 26 ));
FA_296 : FA port map(internal_3_0( 26 ), internal_3_1( 26 ), internal_3_2( 26 ), internal_4_0( 26 ), internal_4_1( 27 ));
FA_297 : FA port map(internal_3_3( 26 ), internal_3_4( 26 ), internal_3_5( 26 ), internal_4_0( 26 ), internal_4_1( 27 ));
FA_298 : FA port map(internal_3_0( 27 ), internal_3_1( 27 ), internal_3_2( 27 ), internal_4_0( 27 ), internal_4_1( 28 ));
FA_299 : FA port map(internal_3_3( 27 ), internal_3_4( 27 ), internal_3_5( 27 ), internal_4_0( 27 ), internal_4_1( 28 ));
FA_300 : FA port map(internal_3_0( 28 ), internal_3_1( 28 ), internal_3_2( 28 ), internal_4_0( 28 ), internal_4_1( 29 ));
FA_301 : FA port map(internal_3_3( 28 ), internal_3_4( 28 ), internal_3_5( 28 ), internal_4_0( 28 ), internal_4_1( 29 ));
FA_302 : FA port map(internal_3_0( 29 ), internal_3_1( 29 ), internal_3_2( 29 ), internal_4_0( 29 ), internal_4_1( 30 ));
FA_303 : FA port map(internal_3_3( 29 ), internal_3_4( 29 ), internal_3_5( 29 ), internal_4_0( 29 ), internal_4_1( 30 ));
FA_304 : FA port map(internal_3_0( 30 ), internal_3_1( 30 ), internal_3_2( 30 ), internal_4_0( 30 ), internal_4_1( 31 ));
FA_305 : FA port map(internal_3_3( 30 ), internal_3_4( 30 ), internal_3_5( 30 ), internal_4_0( 30 ), internal_4_1( 31 ));
FA_306 : FA port map(internal_3_0( 31 ), internal_3_1( 31 ), internal_3_2( 31 ), internal_4_0( 31 ), internal_4_1( 32 ));
FA_307 : FA port map(internal_3_3( 31 ), internal_3_4( 31 ), internal_3_5( 31 ), internal_4_0( 31 ), internal_4_1( 32 ));
FA_308 : FA port map(internal_3_0( 32 ), internal_3_1( 32 ), internal_3_2( 32 ), internal_4_0( 32 ), internal_4_1( 33 ));
FA_309 : FA port map(internal_3_3( 32 ), internal_3_4( 32 ), internal_3_5( 32 ), internal_4_0( 32 ), internal_4_1( 33 ));
FA_310 : FA port map(internal_3_0( 33 ), internal_3_1( 33 ), internal_3_2( 33 ), internal_4_0( 33 ), internal_4_1( 34 ));
FA_311 : FA port map(internal_3_3( 33 ), internal_3_4( 33 ), internal_3_5( 33 ), internal_4_0( 33 ), internal_4_1( 34 ));
FA_312 : FA port map(internal_3_0( 34 ), internal_3_1( 34 ), internal_3_2( 34 ), internal_4_0( 34 ), internal_4_1( 35 ));
FA_313 : FA port map(internal_3_3( 34 ), internal_3_4( 34 ), internal_3_5( 34 ), internal_4_0( 34 ), internal_4_1( 35 ));
FA_314 : FA port map(internal_3_0( 35 ), internal_3_1( 35 ), internal_3_2( 35 ), internal_4_0( 35 ), internal_4_1( 36 ));
FA_315 : FA port map(internal_3_3( 35 ), internal_3_4( 35 ), internal_3_5( 35 ), internal_4_0( 35 ), internal_4_1( 36 ));
FA_316 : FA port map(internal_3_0( 36 ), internal_3_1( 36 ), internal_3_2( 36 ), internal_4_0( 36 ), internal_4_1( 37 ));
FA_317 : FA port map(internal_3_3( 36 ), internal_3_4( 36 ), internal_3_5( 36 ), internal_4_0( 36 ), internal_4_1( 37 ));
FA_318 : FA port map(internal_3_0( 37 ), internal_3_1( 37 ), internal_3_2( 37 ), internal_4_0( 37 ), internal_4_1( 38 ));
FA_319 : FA port map(internal_3_3( 37 ), internal_3_4( 37 ), internal_3_5( 37 ), internal_4_0( 37 ), internal_4_1( 38 ));
FA_320 : FA port map(internal_3_0( 38 ), internal_3_1( 38 ), internal_3_2( 38 ), internal_4_0( 38 ), internal_4_1( 39 ));
FA_321 : FA port map(internal_3_3( 38 ), internal_3_4( 38 ), internal_3_5( 38 ), internal_4_0( 38 ), internal_4_1( 39 ));
FA_322 : FA port map(internal_3_0( 39 ), internal_3_1( 39 ), internal_3_2( 39 ), internal_4_0( 39 ), internal_4_1( 40 ));
FA_323 : FA port map(internal_3_3( 39 ), internal_3_4( 39 ), internal_3_5( 39 ), internal_4_0( 39 ), internal_4_1( 40 ));
FA_324 : FA port map(internal_3_0( 40 ), internal_3_1( 40 ), internal_3_2( 40 ), internal_4_0( 40 ), internal_4_1( 41 ));
FA_325 : FA port map(internal_3_3( 40 ), internal_3_4( 40 ), internal_3_5( 40 ), internal_4_0( 40 ), internal_4_1( 41 ));
FA_326 : FA port map(internal_3_0( 41 ), internal_3_1( 41 ), internal_3_2( 41 ), internal_4_0( 41 ), internal_4_1( 42 ));
FA_327 : FA port map(internal_3_3( 41 ), internal_3_4( 41 ), internal_3_5( 41 ), internal_4_0( 41 ), internal_4_1( 42 ));
FA_328 : FA port map(internal_3_0( 42 ), internal_3_1( 42 ), internal_3_2( 42 ), internal_4_0( 42 ), internal_4_1( 43 ));
FA_329 : FA port map(internal_3_3( 42 ), internal_3_4( 42 ), internal_3_5( 42 ), internal_4_0( 42 ), internal_4_1( 43 ));
FA_330 : FA port map(internal_3_0( 43 ), internal_3_1( 43 ), internal_3_2( 43 ), internal_4_0( 43 ), internal_4_1( 44 ));
FA_331 : FA port map(internal_3_3( 43 ), internal_3_4( 43 ), internal_3_5( 43 ), internal_4_0( 43 ), internal_4_1( 44 ));
FA_332 : FA port map(internal_3_0( 44 ), internal_3_1( 44 ), internal_3_2( 44 ), internal_4_0( 44 ), internal_4_1( 45 ));
FA_333 : FA port map(internal_3_3( 44 ), internal_3_4( 44 ), internal_3_5( 44 ), internal_4_0( 44 ), internal_4_1( 45 ));
FA_334 : FA port map(internal_3_0( 45 ), internal_3_1( 45 ), internal_3_2( 45 ), internal_4_0( 45 ), internal_4_1( 46 ));
FA_335 : FA port map(internal_3_3( 45 ), internal_3_4( 45 ), internal_3_5( 45 ), internal_4_0( 45 ), internal_4_1( 46 ));
FA_336 : FA port map(internal_3_0( 46 ), internal_3_1( 46 ), internal_3_2( 46 ), internal_4_0( 46 ), internal_4_1( 47 ));
FA_337 : FA port map(internal_3_3( 46 ), internal_3_4( 46 ), internal_3_5( 46 ), internal_4_0( 46 ), internal_4_1( 47 ));
FA_338 : FA port map(internal_3_0( 47 ), internal_3_1( 47 ), internal_3_2( 47 ), internal_4_0( 47 ), internal_4_1( 48 ));
FA_339 : FA port map(internal_3_3( 47 ), internal_3_4( 47 ), internal_3_5( 47 ), internal_4_0( 47 ), internal_4_1( 48 ));
FA_340 : FA port map(internal_3_0( 48 ), internal_3_1( 48 ), internal_3_2( 48 ), internal_4_0( 48 ), internal_4_1( 49 ));
FA_341 : FA port map(internal_3_3( 48 ), internal_3_4( 48 ), internal_3_5( 48 ), internal_4_0( 48 ), internal_4_1( 49 ));
FA_342 : FA port map(internal_3_0( 49 ), internal_3_1( 49 ), internal_3_2( 49 ), internal_4_0( 49 ), internal_4_1( 50 ));
FA_343 : FA port map(internal_3_3( 49 ), internal_3_4( 49 ), internal_3_5( 49 ), internal_4_0( 49 ), internal_4_1( 50 ));
FA_344 : FA port map(internal_3_0( 50 ), internal_3_1( 50 ), internal_3_2( 50 ), internal_4_0( 50 ), internal_4_1( 51 ));
FA_345 : FA port map(internal_3_3( 50 ), internal_3_4( 50 ), internal_3_5( 50 ), internal_4_0( 50 ), internal_4_1( 51 ));
FA_346 : FA port map(internal_3_0( 51 ), internal_3_1( 51 ), internal_3_2( 51 ), internal_4_0( 51 ), internal_4_1( 52 ));
FA_347 : FA port map(internal_3_3( 51 ), internal_3_4( 51 ), internal_3_5( 51 ), internal_4_0( 51 ), internal_4_1( 52 ));
FA_348 : FA port map(internal_3_0( 52 ), internal_3_1( 52 ), internal_3_2( 52 ), internal_4_0( 52 ), internal_4_1( 53 ));
FA_349 : FA port map(internal_3_3( 52 ), internal_3_4( 52 ), internal_3_5( 52 ), internal_4_0( 52 ), internal_4_1( 53 ));
FA_350 : FA port map(internal_3_0( 53 ), internal_3_1( 53 ), internal_3_2( 53 ), internal_4_0( 53 ), internal_4_1( 54 ));
FA_351 : FA port map(internal_3_3( 53 ), internal_3_4( 53 ), internal_3_5( 53 ), internal_4_0( 53 ), internal_4_1( 54 ));
FA_352 : FA port map(internal_3_0( 54 ), internal_3_1( 54 ), internal_3_2( 54 ), internal_4_0( 54 ), internal_4_1( 55 ));
FA_353 : FA port map(internal_3_3( 54 ), internal_3_4( 54 ), internal_3_5( 54 ), internal_4_0( 54 ), internal_4_1( 55 ));
FA_354 : FA port map(internal_3_0( 55 ), internal_3_1( 55 ), internal_3_2( 55 ), internal_4_0( 55 ), internal_4_1( 56 ));
FA_355 : FA port map(internal_3_3( 55 ), internal_3_4( 55 ), internal_3_5( 55 ), internal_4_0( 55 ), internal_4_1( 56 ));
FA_356 : FA port map(internal_3_0( 56 ), internal_3_1( 56 ), internal_3_2( 56 ), internal_4_0( 56 ), internal_4_1( 57 ));
FA_357 : FA port map(internal_3_3( 56 ), internal_3_4( 56 ), internal_3_5( 56 ), internal_4_0( 56 ), internal_4_1( 57 ));
FA_358 : FA port map(internal_3_0( 57 ), internal_3_1( 57 ), internal_3_2( 57 ), internal_4_0( 57 ), internal_4_1( 58 ));
HA_39 : HA port map(internal_3_3( 57 ), internal_3_4( 57 ), internal_4_1( 57 ), internal_4_2( 58 ));
FA_359 : FA port map(internal_3_0( 58 ), internal_3_1( 58 ), internal_3_2( 58 ), internal_4_0( 58 ), internal_4_1( 59 ));
HA_40 : HA port map(internal_3_3( 58 ), internal_3_4( 58 ), internal_4_1( 58 ), internal_4_2( 59 ));
FA_360 : FA port map(internal_3_0( 59 ), internal_3_1( 59 ), internal_3_2( 59 ), internal_4_0( 59 ), internal_4_1( 60 ));
HA_41 : HA port map(internal_3_0( 60 ), internal_3_1( 60 ), internal_4_0( 60 ), internal_4_1( 61 ));
HA_42 : HA port map(internal_4_0( 4 ), internal_4_1( 4 ), internal_5_0( 4 ), internal_5_1( 5 ));
HA_43 : HA port map(internal_4_0( 5 ), internal_4_1( 5 ), internal_5_0( 5 ), internal_5_1( 6 ));
FA_361 : FA port map(internal_4_0( 6 ), internal_4_1( 6 ), internal_4_2( 6 ), internal_5_0( 6 ), internal_5_1( 7 ));
FA_362 : FA port map(internal_4_0( 7 ), internal_4_1( 7 ), internal_4_2( 7 ), internal_5_0( 7 ), internal_5_1( 8 ));
FA_363 : FA port map(internal_4_0( 8 ), internal_4_1( 8 ), internal_4_2( 8 ), internal_5_0( 8 ), internal_5_1( 9 ));
FA_364 : FA port map(internal_4_0( 9 ), internal_4_1( 9 ), internal_4_2( 9 ), internal_5_0( 9 ), internal_5_1( 10 ));
FA_365 : FA port map(internal_4_0( 10 ), internal_4_1( 10 ), internal_4_2( 10 ), internal_5_0( 10 ), internal_5_1( 11 ));
FA_366 : FA port map(internal_4_0( 11 ), internal_4_1( 11 ), internal_4_2( 11 ), internal_5_0( 11 ), internal_5_1( 12 ));
FA_367 : FA port map(internal_4_0( 12 ), internal_4_1( 12 ), internal_4_2( 12 ), internal_5_0( 12 ), internal_5_1( 13 ));
FA_368 : FA port map(internal_4_0( 13 ), internal_4_1( 13 ), internal_4_2( 13 ), internal_5_0( 13 ), internal_5_1( 14 ));
FA_369 : FA port map(internal_4_0( 14 ), internal_4_1( 14 ), internal_4_2( 14 ), internal_5_0( 14 ), internal_5_1( 15 ));
FA_370 : FA port map(internal_4_0( 15 ), internal_4_1( 15 ), internal_4_2( 15 ), internal_5_0( 15 ), internal_5_1( 16 ));
FA_371 : FA port map(internal_4_0( 16 ), internal_4_1( 16 ), internal_4_2( 16 ), internal_5_0( 16 ), internal_5_1( 17 ));
FA_372 : FA port map(internal_4_0( 17 ), internal_4_1( 17 ), internal_4_2( 17 ), internal_5_0( 17 ), internal_5_1( 18 ));
FA_373 : FA port map(internal_4_0( 18 ), internal_4_1( 18 ), internal_4_2( 18 ), internal_5_0( 18 ), internal_5_1( 19 ));
FA_374 : FA port map(internal_4_0( 19 ), internal_4_1( 19 ), internal_4_2( 19 ), internal_5_0( 19 ), internal_5_1( 20 ));
FA_375 : FA port map(internal_4_0( 20 ), internal_4_1( 20 ), internal_4_2( 20 ), internal_5_0( 20 ), internal_5_1( 21 ));
FA_376 : FA port map(internal_4_0( 21 ), internal_4_1( 21 ), internal_4_2( 21 ), internal_5_0( 21 ), internal_5_1( 22 ));
FA_377 : FA port map(internal_4_0( 22 ), internal_4_1( 22 ), internal_4_2( 22 ), internal_5_0( 22 ), internal_5_1( 23 ));
FA_378 : FA port map(internal_4_0( 23 ), internal_4_1( 23 ), internal_4_2( 23 ), internal_5_0( 23 ), internal_5_1( 24 ));
FA_379 : FA port map(internal_4_0( 24 ), internal_4_1( 24 ), internal_4_2( 24 ), internal_5_0( 24 ), internal_5_1( 25 ));
FA_380 : FA port map(internal_4_0( 25 ), internal_4_1( 25 ), internal_4_2( 25 ), internal_5_0( 25 ), internal_5_1( 26 ));
FA_381 : FA port map(internal_4_0( 26 ), internal_4_1( 26 ), internal_4_2( 26 ), internal_5_0( 26 ), internal_5_1( 27 ));
FA_382 : FA port map(internal_4_0( 27 ), internal_4_1( 27 ), internal_4_2( 27 ), internal_5_0( 27 ), internal_5_1( 28 ));
FA_383 : FA port map(internal_4_0( 28 ), internal_4_1( 28 ), internal_4_2( 28 ), internal_5_0( 28 ), internal_5_1( 29 ));
FA_384 : FA port map(internal_4_0( 29 ), internal_4_1( 29 ), internal_4_2( 29 ), internal_5_0( 29 ), internal_5_1( 30 ));
FA_385 : FA port map(internal_4_0( 30 ), internal_4_1( 30 ), internal_4_2( 30 ), internal_5_0( 30 ), internal_5_1( 31 ));
FA_386 : FA port map(internal_4_0( 31 ), internal_4_1( 31 ), internal_4_2( 31 ), internal_5_0( 31 ), internal_5_1( 32 ));
FA_387 : FA port map(internal_4_0( 32 ), internal_4_1( 32 ), internal_4_2( 32 ), internal_5_0( 32 ), internal_5_1( 33 ));
FA_388 : FA port map(internal_4_0( 33 ), internal_4_1( 33 ), internal_4_2( 33 ), internal_5_0( 33 ), internal_5_1( 34 ));
FA_389 : FA port map(internal_4_0( 34 ), internal_4_1( 34 ), internal_4_2( 34 ), internal_5_0( 34 ), internal_5_1( 35 ));
FA_390 : FA port map(internal_4_0( 35 ), internal_4_1( 35 ), internal_4_2( 35 ), internal_5_0( 35 ), internal_5_1( 36 ));
FA_391 : FA port map(internal_4_0( 36 ), internal_4_1( 36 ), internal_4_2( 36 ), internal_5_0( 36 ), internal_5_1( 37 ));
FA_392 : FA port map(internal_4_0( 37 ), internal_4_1( 37 ), internal_4_2( 37 ), internal_5_0( 37 ), internal_5_1( 38 ));
FA_393 : FA port map(internal_4_0( 38 ), internal_4_1( 38 ), internal_4_2( 38 ), internal_5_0( 38 ), internal_5_1( 39 ));
FA_394 : FA port map(internal_4_0( 39 ), internal_4_1( 39 ), internal_4_2( 39 ), internal_5_0( 39 ), internal_5_1( 40 ));
FA_395 : FA port map(internal_4_0( 40 ), internal_4_1( 40 ), internal_4_2( 40 ), internal_5_0( 40 ), internal_5_1( 41 ));
FA_396 : FA port map(internal_4_0( 41 ), internal_4_1( 41 ), internal_4_2( 41 ), internal_5_0( 41 ), internal_5_1( 42 ));
FA_397 : FA port map(internal_4_0( 42 ), internal_4_1( 42 ), internal_4_2( 42 ), internal_5_0( 42 ), internal_5_1( 43 ));
FA_398 : FA port map(internal_4_0( 43 ), internal_4_1( 43 ), internal_4_2( 43 ), internal_5_0( 43 ), internal_5_1( 44 ));
FA_399 : FA port map(internal_4_0( 44 ), internal_4_1( 44 ), internal_4_2( 44 ), internal_5_0( 44 ), internal_5_1( 45 ));
FA_400 : FA port map(internal_4_0( 45 ), internal_4_1( 45 ), internal_4_2( 45 ), internal_5_0( 45 ), internal_5_1( 46 ));
FA_401 : FA port map(internal_4_0( 46 ), internal_4_1( 46 ), internal_4_2( 46 ), internal_5_0( 46 ), internal_5_1( 47 ));
FA_402 : FA port map(internal_4_0( 47 ), internal_4_1( 47 ), internal_4_2( 47 ), internal_5_0( 47 ), internal_5_1( 48 ));
FA_403 : FA port map(internal_4_0( 48 ), internal_4_1( 48 ), internal_4_2( 48 ), internal_5_0( 48 ), internal_5_1( 49 ));
FA_404 : FA port map(internal_4_0( 49 ), internal_4_1( 49 ), internal_4_2( 49 ), internal_5_0( 49 ), internal_5_1( 50 ));
FA_405 : FA port map(internal_4_0( 50 ), internal_4_1( 50 ), internal_4_2( 50 ), internal_5_0( 50 ), internal_5_1( 51 ));
FA_406 : FA port map(internal_4_0( 51 ), internal_4_1( 51 ), internal_4_2( 51 ), internal_5_0( 51 ), internal_5_1( 52 ));
FA_407 : FA port map(internal_4_0( 52 ), internal_4_1( 52 ), internal_4_2( 52 ), internal_5_0( 52 ), internal_5_1( 53 ));
FA_408 : FA port map(internal_4_0( 53 ), internal_4_1( 53 ), internal_4_2( 53 ), internal_5_0( 53 ), internal_5_1( 54 ));
FA_409 : FA port map(internal_4_0( 54 ), internal_4_1( 54 ), internal_4_2( 54 ), internal_5_0( 54 ), internal_5_1( 55 ));
FA_410 : FA port map(internal_4_0( 55 ), internal_4_1( 55 ), internal_4_2( 55 ), internal_5_0( 55 ), internal_5_1( 56 ));
FA_411 : FA port map(internal_4_0( 56 ), internal_4_1( 56 ), internal_4_2( 56 ), internal_5_0( 56 ), internal_5_1( 57 ));
FA_412 : FA port map(internal_4_0( 57 ), internal_4_1( 57 ), internal_4_2( 57 ), internal_5_0( 57 ), internal_5_1( 58 ));
FA_413 : FA port map(internal_4_0( 58 ), internal_4_1( 58 ), internal_4_2( 58 ), internal_5_0( 58 ), internal_5_1( 59 ));
FA_414 : FA port map(internal_4_0( 59 ), internal_4_1( 59 ), internal_4_2( 59 ), internal_5_0( 59 ), internal_5_1( 60 ));
FA_415 : FA port map(internal_4_0( 60 ), internal_4_1( 60 ), internal_4_2( 60 ), internal_5_0( 60 ), internal_5_1( 61 ));
HA_44 : HA port map(internal_4_0( 61 ), internal_4_1( 61 ), internal_5_0( 61 ), internal_5_1( 62 ));
HA_45 : HA port map(internal_4_0( 62 ), internal_4_1( 62 ), internal_5_0( 62 ), internal_5_1( 63 ));
HA_46 : HA port map(internal_5_0( 2 ), internal_5_1( 2 ), internal_6_0( 2 ), internal_6_1( 3 ));
HA_47 : HA port map(internal_5_0( 3 ), internal_5_1( 3 ), internal_6_0( 3 ), internal_6_1( 4 ));
FA_416 : FA port map(internal_5_0( 4 ), internal_5_1( 4 ), internal_5_2( 4 ), internal_6_0( 4 ), internal_6_1( 5 ));
FA_417 : FA port map(internal_5_0( 5 ), internal_5_1( 5 ), internal_5_2( 5 ), internal_6_0( 5 ), internal_6_1( 6 ));
FA_418 : FA port map(internal_5_0( 6 ), internal_5_1( 6 ), internal_5_2( 6 ), internal_6_0( 6 ), internal_6_1( 7 ));
FA_419 : FA port map(internal_5_0( 7 ), internal_5_1( 7 ), internal_5_2( 7 ), internal_6_0( 7 ), internal_6_1( 8 ));
FA_420 : FA port map(internal_5_0( 8 ), internal_5_1( 8 ), internal_5_2( 8 ), internal_6_0( 8 ), internal_6_1( 9 ));
FA_421 : FA port map(internal_5_0( 9 ), internal_5_1( 9 ), internal_5_2( 9 ), internal_6_0( 9 ), internal_6_1( 10 ));
FA_422 : FA port map(internal_5_0( 10 ), internal_5_1( 10 ), internal_5_2( 10 ), internal_6_0( 10 ), internal_6_1( 11 ));
FA_423 : FA port map(internal_5_0( 11 ), internal_5_1( 11 ), internal_5_2( 11 ), internal_6_0( 11 ), internal_6_1( 12 ));
FA_424 : FA port map(internal_5_0( 12 ), internal_5_1( 12 ), internal_5_2( 12 ), internal_6_0( 12 ), internal_6_1( 13 ));
FA_425 : FA port map(internal_5_0( 13 ), internal_5_1( 13 ), internal_5_2( 13 ), internal_6_0( 13 ), internal_6_1( 14 ));
FA_426 : FA port map(internal_5_0( 14 ), internal_5_1( 14 ), internal_5_2( 14 ), internal_6_0( 14 ), internal_6_1( 15 ));
FA_427 : FA port map(internal_5_0( 15 ), internal_5_1( 15 ), internal_5_2( 15 ), internal_6_0( 15 ), internal_6_1( 16 ));
FA_428 : FA port map(internal_5_0( 16 ), internal_5_1( 16 ), internal_5_2( 16 ), internal_6_0( 16 ), internal_6_1( 17 ));
FA_429 : FA port map(internal_5_0( 17 ), internal_5_1( 17 ), internal_5_2( 17 ), internal_6_0( 17 ), internal_6_1( 18 ));
FA_430 : FA port map(internal_5_0( 18 ), internal_5_1( 18 ), internal_5_2( 18 ), internal_6_0( 18 ), internal_6_1( 19 ));
FA_431 : FA port map(internal_5_0( 19 ), internal_5_1( 19 ), internal_5_2( 19 ), internal_6_0( 19 ), internal_6_1( 20 ));
FA_432 : FA port map(internal_5_0( 20 ), internal_5_1( 20 ), internal_5_2( 20 ), internal_6_0( 20 ), internal_6_1( 21 ));
FA_433 : FA port map(internal_5_0( 21 ), internal_5_1( 21 ), internal_5_2( 21 ), internal_6_0( 21 ), internal_6_1( 22 ));
FA_434 : FA port map(internal_5_0( 22 ), internal_5_1( 22 ), internal_5_2( 22 ), internal_6_0( 22 ), internal_6_1( 23 ));
FA_435 : FA port map(internal_5_0( 23 ), internal_5_1( 23 ), internal_5_2( 23 ), internal_6_0( 23 ), internal_6_1( 24 ));
FA_436 : FA port map(internal_5_0( 24 ), internal_5_1( 24 ), internal_5_2( 24 ), internal_6_0( 24 ), internal_6_1( 25 ));
FA_437 : FA port map(internal_5_0( 25 ), internal_5_1( 25 ), internal_5_2( 25 ), internal_6_0( 25 ), internal_6_1( 26 ));
FA_438 : FA port map(internal_5_0( 26 ), internal_5_1( 26 ), internal_5_2( 26 ), internal_6_0( 26 ), internal_6_1( 27 ));
FA_439 : FA port map(internal_5_0( 27 ), internal_5_1( 27 ), internal_5_2( 27 ), internal_6_0( 27 ), internal_6_1( 28 ));
FA_440 : FA port map(internal_5_0( 28 ), internal_5_1( 28 ), internal_5_2( 28 ), internal_6_0( 28 ), internal_6_1( 29 ));
FA_441 : FA port map(internal_5_0( 29 ), internal_5_1( 29 ), internal_5_2( 29 ), internal_6_0( 29 ), internal_6_1( 30 ));
FA_442 : FA port map(internal_5_0( 30 ), internal_5_1( 30 ), internal_5_2( 30 ), internal_6_0( 30 ), internal_6_1( 31 ));
FA_443 : FA port map(internal_5_0( 31 ), internal_5_1( 31 ), internal_5_2( 31 ), internal_6_0( 31 ), internal_6_1( 32 ));
FA_444 : FA port map(internal_5_0( 32 ), internal_5_1( 32 ), internal_5_2( 32 ), internal_6_0( 32 ), internal_6_1( 33 ));
FA_445 : FA port map(internal_5_0( 33 ), internal_5_1( 33 ), internal_5_2( 33 ), internal_6_0( 33 ), internal_6_1( 34 ));
FA_446 : FA port map(internal_5_0( 34 ), internal_5_1( 34 ), internal_5_2( 34 ), internal_6_0( 34 ), internal_6_1( 35 ));
FA_447 : FA port map(internal_5_0( 35 ), internal_5_1( 35 ), internal_5_2( 35 ), internal_6_0( 35 ), internal_6_1( 36 ));
FA_448 : FA port map(internal_5_0( 36 ), internal_5_1( 36 ), internal_5_2( 36 ), internal_6_0( 36 ), internal_6_1( 37 ));
FA_449 : FA port map(internal_5_0( 37 ), internal_5_1( 37 ), internal_5_2( 37 ), internal_6_0( 37 ), internal_6_1( 38 ));
FA_450 : FA port map(internal_5_0( 38 ), internal_5_1( 38 ), internal_5_2( 38 ), internal_6_0( 38 ), internal_6_1( 39 ));
FA_451 : FA port map(internal_5_0( 39 ), internal_5_1( 39 ), internal_5_2( 39 ), internal_6_0( 39 ), internal_6_1( 40 ));
FA_452 : FA port map(internal_5_0( 40 ), internal_5_1( 40 ), internal_5_2( 40 ), internal_6_0( 40 ), internal_6_1( 41 ));
FA_453 : FA port map(internal_5_0( 41 ), internal_5_1( 41 ), internal_5_2( 41 ), internal_6_0( 41 ), internal_6_1( 42 ));
FA_454 : FA port map(internal_5_0( 42 ), internal_5_1( 42 ), internal_5_2( 42 ), internal_6_0( 42 ), internal_6_1( 43 ));
FA_455 : FA port map(internal_5_0( 43 ), internal_5_1( 43 ), internal_5_2( 43 ), internal_6_0( 43 ), internal_6_1( 44 ));
FA_456 : FA port map(internal_5_0( 44 ), internal_5_1( 44 ), internal_5_2( 44 ), internal_6_0( 44 ), internal_6_1( 45 ));
FA_457 : FA port map(internal_5_0( 45 ), internal_5_1( 45 ), internal_5_2( 45 ), internal_6_0( 45 ), internal_6_1( 46 ));
FA_458 : FA port map(internal_5_0( 46 ), internal_5_1( 46 ), internal_5_2( 46 ), internal_6_0( 46 ), internal_6_1( 47 ));
FA_459 : FA port map(internal_5_0( 47 ), internal_5_1( 47 ), internal_5_2( 47 ), internal_6_0( 47 ), internal_6_1( 48 ));
FA_460 : FA port map(internal_5_0( 48 ), internal_5_1( 48 ), internal_5_2( 48 ), internal_6_0( 48 ), internal_6_1( 49 ));
FA_461 : FA port map(internal_5_0( 49 ), internal_5_1( 49 ), internal_5_2( 49 ), internal_6_0( 49 ), internal_6_1( 50 ));
FA_462 : FA port map(internal_5_0( 50 ), internal_5_1( 50 ), internal_5_2( 50 ), internal_6_0( 50 ), internal_6_1( 51 ));
FA_463 : FA port map(internal_5_0( 51 ), internal_5_1( 51 ), internal_5_2( 51 ), internal_6_0( 51 ), internal_6_1( 52 ));
FA_464 : FA port map(internal_5_0( 52 ), internal_5_1( 52 ), internal_5_2( 52 ), internal_6_0( 52 ), internal_6_1( 53 ));
FA_465 : FA port map(internal_5_0( 53 ), internal_5_1( 53 ), internal_5_2( 53 ), internal_6_0( 53 ), internal_6_1( 54 ));
FA_466 : FA port map(internal_5_0( 54 ), internal_5_1( 54 ), internal_5_2( 54 ), internal_6_0( 54 ), internal_6_1( 55 ));
FA_467 : FA port map(internal_5_0( 55 ), internal_5_1( 55 ), internal_5_2( 55 ), internal_6_0( 55 ), internal_6_1( 56 ));
FA_468 : FA port map(internal_5_0( 56 ), internal_5_1( 56 ), internal_5_2( 56 ), internal_6_0( 56 ), internal_6_1( 57 ));
FA_469 : FA port map(internal_5_0( 57 ), internal_5_1( 57 ), internal_5_2( 57 ), internal_6_0( 57 ), internal_6_1( 58 ));
FA_470 : FA port map(internal_5_0( 58 ), internal_5_1( 58 ), internal_5_2( 58 ), internal_6_0( 58 ), internal_6_1( 59 ));
FA_471 : FA port map(internal_5_0( 59 ), internal_5_1( 59 ), internal_5_2( 59 ), internal_6_0( 59 ), internal_6_1( 60 ));
FA_472 : FA port map(internal_5_0( 60 ), internal_5_1( 60 ), internal_5_2( 60 ), internal_6_0( 60 ), internal_6_1( 61 ));
FA_473 : FA port map(internal_5_0( 61 ), internal_5_1( 61 ), internal_5_2( 61 ), internal_6_0( 61 ), internal_6_1( 62 ));
FA_474 : FA port map(internal_5_0( 62 ), internal_5_1( 62 ), internal_5_2( 62 ), internal_6_0( 62 ), internal_6_1( 63 ));
HA_48 : HA port map(internal_5_0( 63 ), internal_5_1( 63 ), internal_6_0( 63 ), internal_6_1( 64 ));


end architecture ;