LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY FA IS
PORT(
		A, B, Cin : IN STD_LOGIC;
		S, Co : OUT STD_LOGIC
	 );	
END FULL_ADDER;

ARCHITECTURE structural OF FULL_ADDER IS

SIGNAL OUT_FIRST_1, OUT_FIRST_2, OUT_SECOND : STD_LOGIC;

	COMPONENT HA 
	PORT(
		A, B : IN STD_LOGIC;
		SUM, CARRY : OUT STD_LOGIC
	 );
	END COMPONENT;
	
BEGIN

HALF1 : HA PORT MAP (IN_1 => A, IN_2 => B, CARRY => OUT_FIRST_2, SUM => OUT_FIRST_1);
HALF2 : HA PORT MAP (IN_1 => Cin, IN_2 => OUT_FIRST_1, CARRY => OUT_SECOND, SUM => S);
Co <= OUT_SECOND OR OUT_FIRST_2;

END BEHAVIOUR;
	