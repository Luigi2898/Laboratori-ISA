LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY REG IS
	PORT(REG_IN : IN signed(10 DOWNTO 0);
		 REG_OUT : OUT signed(10 DOWNTO 0);
		 CLK, RST_N, LOAD : IN STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEH OF REG IS

BEGIN
REGPROC: PROCESS(CLK, RST_N)
BEGIN
IF(RST_N = '0') THEN
	REG_OUT <= (OTHERS => '0');
     ELSIF(CLK'EVENT AND CLK = '1') THEN
		 IF(LOAD = '1') THEN
		 REG_OUT <= REG_IN;
		 END IF;
END IF;

END PROCESS;

END ARCHITECTURE;
