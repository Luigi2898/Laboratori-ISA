`timescale 10 ns/ 1 ns

module tb_HDU();

	reg ID_EX_MEMREAD_IN = 1'b0;
	reg [31:0] INSTR_IF_ID_IN = 32'b11111111110000010000000100010011;
    reg [31:0] INSTR_ID_EX_IN = 32'b00000000101000000000001010010011;
    wire IF_ID_EN_OUT;
	wire PC_EN_OUT;
	wire CTRL_BUBBLE_OUT;

    HDU     DUT(.INSTR_IF_ID_IN(INSTR_IF_ID_IN),
                .INSTR_ID_EX_IN(INSTR_ID_EX_IN),
                .ID_EX_MEMREAD_IN(ID_EX_MEMREAD_IN),
                .IF_ID_EN_OUT(IF_ID_EN_OUT),
                .PC_EN_OUT(PC_EN_OUT),
                .CTRL_BUBBLE_OUT(CTRL_BUBBLE_OUT));
    initial 
    begin 
	#10 ID_EX_MEMREAD_IN = 1'b0;
        INSTR_IF_ID_IN = 32'b00000000010100010010000000100011;
        INSTR_ID_EX_IN = 32'b11111111110000010000000100010011;
	#20 ID_EX_MEMREAD_IN = 1'b0;
        INSTR_IF_ID_IN = 32'b00000000010100101000001100110011;
        INSTR_ID_EX_IN = 32'b00000000010100010010000000100011;
    #30 ID_EX_MEMREAD_IN = 1'b0;
        INSTR_IF_ID_IN = 32'b00000000000000010010001010000011;
        INSTR_ID_EX_IN = 32'b00000000010100101000001100110011; 
    #40 ID_EX_MEMREAD_IN = 1'b1;
        INSTR_IF_ID_IN = 32'b00000000000000101000001100110011;
        INSTR_ID_EX_IN = 32'b00000000000000010010001010000011;
    #50 ID_EX_MEMREAD_IN = 1'b1;
        INSTR_IF_ID_IN = 32'b00000000000000000000001100110011;
        INSTR_ID_EX_IN = 32'b00000000000000010010001010000011;            
	end
            

    
endmodule
