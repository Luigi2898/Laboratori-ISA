library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity ALU is
  port (
  
  );
end entity;

architecture arch of ALU is

begin

end architecture;
