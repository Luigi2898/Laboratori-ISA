library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity BPU is
  port (
    clock : in std_logic
  );
end entity;

architecture arch of BPU is

begin

end architecture;
