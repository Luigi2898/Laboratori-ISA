LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY HA IS
PORT(
		A, B : IN STD_LOGIC;
		SUM, CARRY : OUT STD_LOGIC
	 );
END HA;

ARCHITECTURE struct OF HA IS
BEGIN
SUM <= A XOR B;
CARRY <= A AND B;
END BEHAVIOUR;