module mult(   input logic [31:0] A, B, 
                output logic [31:0] OUT );

    assign OUT = A * B;

endmodule: mult
