library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity HDU is
  port (
    clock : in std_logic
  );
end entity;

architecture arch of HDU is

begin

end architecture;
