library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity DADDA is
  port (
    
  ) ;
end DADDA ; 

architecture structural of DADDA is

begin

end architecture ;