library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity CU is
  port (
    OPCODE : in std_logic_vector(6 downto 0)
  );
end entity;

architecture arch of CU is

begin

end architecture;
