library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity CU is
  port (
    clock : in std_logic
  );
end entity;

architecture arch of CU is

begin

end architecture;
